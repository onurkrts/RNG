magic
tech sky130A
magscale 1 2
timestamp 1647847231
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 283834 700748 283840 700800
rect 283892 700788 283898 700800
rect 328454 700788 328460 700800
rect 283892 700760 328460 700788
rect 283892 700748 283898 700760
rect 328454 700748 328460 700760
rect 328512 700748 328518 700800
rect 318794 700680 318800 700732
rect 318852 700720 318858 700732
rect 413646 700720 413652 700732
rect 318852 700692 413652 700720
rect 318852 700680 318858 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 218974 700612 218980 700664
rect 219032 700652 219038 700664
rect 332594 700652 332600 700664
rect 219032 700624 332600 700652
rect 219032 700612 219038 700624
rect 332594 700612 332600 700624
rect 332652 700612 332658 700664
rect 154114 700544 154120 700596
rect 154172 700584 154178 700596
rect 338114 700584 338120 700596
rect 154172 700556 338120 700584
rect 154172 700544 154178 700556
rect 338114 700544 338120 700556
rect 338172 700544 338178 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 342254 700516 342260 700528
rect 89220 700488 342260 700516
rect 89220 700476 89226 700488
rect 342254 700476 342260 700488
rect 342312 700476 342318 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 340874 700448 340880 700460
rect 73028 700420 340880 700448
rect 73028 700408 73034 700420
rect 340874 700408 340880 700420
rect 340932 700408 340938 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 347866 700380 347872 700392
rect 24360 700352 347872 700380
rect 24360 700340 24366 700352
rect 347866 700340 347872 700352
rect 347924 700340 347930 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 460198 700272 460204 700324
rect 460256 700312 460262 700324
rect 559650 700312 559656 700324
rect 460256 700284 559656 700312
rect 460256 700272 460262 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 235166 698912 235172 698964
rect 235224 698952 235230 698964
rect 329834 698952 329840 698964
rect 235224 698924 329840 698952
rect 235224 698912 235230 698924
rect 329834 698912 329840 698924
rect 329892 698912 329898 698964
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 303614 696940 303620 696992
rect 303672 696980 303678 696992
rect 580166 696980 580172 696992
rect 303672 696952 580172 696980
rect 303672 696940 303678 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 304994 683136 305000 683188
rect 305052 683176 305058 683188
rect 580166 683176 580172 683188
rect 305052 683148 580172 683176
rect 305052 683136 305058 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 300854 670760 300860 670812
rect 300912 670800 300918 670812
rect 580166 670800 580172 670812
rect 300912 670772 580172 670800
rect 300912 670760 300918 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 351914 670732 351920 670744
rect 3568 670704 351920 670732
rect 3568 670692 3574 670704
rect 351914 670692 351920 670704
rect 351972 670692 351978 670744
rect 306374 660288 306380 660340
rect 306432 660328 306438 660340
rect 460198 660328 460204 660340
rect 306432 660300 460204 660328
rect 306432 660288 306438 660300
rect 460198 660288 460204 660300
rect 460256 660288 460262 660340
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 350534 656928 350540 656940
rect 3568 656900 350540 656928
rect 3568 656888 3574 656900
rect 350534 656888 350540 656900
rect 350592 656888 350598 656940
rect 298094 643084 298100 643136
rect 298152 643124 298158 643136
rect 580166 643124 580172 643136
rect 298152 643096 580172 643124
rect 298152 643084 298158 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 580166 630680 580172 630692
rect 299624 630652 580172 630680
rect 299624 630640 299630 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3326 618264 3332 618316
rect 3384 618304 3390 618316
rect 356054 618304 356060 618316
rect 3384 618276 356060 618304
rect 3384 618264 3390 618276
rect 356054 618264 356060 618276
rect 356112 618264 356118 618316
rect 296714 616836 296720 616888
rect 296772 616876 296778 616888
rect 580166 616876 580172 616888
rect 296772 616848 580172 616876
rect 296772 616836 296778 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 354674 605860 354680 605872
rect 3384 605832 354680 605860
rect 3384 605820 3390 605832
rect 354674 605820 354680 605832
rect 354732 605820 354738 605872
rect 293954 590656 293960 590708
rect 294012 590696 294018 590708
rect 579798 590696 579804 590708
rect 294012 590668 579804 590696
rect 294012 590656 294018 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 295334 576852 295340 576904
rect 295392 576892 295398 576904
rect 580166 576892 580172 576904
rect 295392 576864 580172 576892
rect 295392 576852 295398 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 361574 565876 361580 565888
rect 3108 565848 361580 565876
rect 3108 565836 3114 565848
rect 361574 565836 361580 565848
rect 361632 565836 361638 565888
rect 292574 563048 292580 563100
rect 292632 563088 292638 563100
rect 579798 563088 579804 563100
rect 292632 563060 579804 563088
rect 292632 563048 292638 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 360194 553432 360200 553444
rect 3384 553404 360200 553432
rect 3384 553392 3390 553404
rect 360194 553392 360200 553404
rect 360252 553392 360258 553444
rect 288434 536800 288440 536852
rect 288492 536840 288498 536852
rect 580166 536840 580172 536852
rect 288492 536812 580172 536840
rect 288492 536800 288498 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 320174 527824 320180 527876
rect 320232 527864 320238 527876
rect 364334 527864 364340 527876
rect 320232 527836 364340 527864
rect 320232 527824 320238 527836
rect 364334 527824 364340 527836
rect 364392 527824 364398 527876
rect 289814 524424 289820 524476
rect 289872 524464 289878 524476
rect 580166 524464 580172 524476
rect 289872 524436 580172 524464
rect 289872 524424 289878 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 365714 514808 365720 514820
rect 3384 514780 365720 514808
rect 3384 514768 3390 514780
rect 365714 514768 365720 514780
rect 365772 514768 365778 514820
rect 287054 510620 287060 510672
rect 287112 510660 287118 510672
rect 580166 510660 580172 510672
rect 287112 510632 580172 510660
rect 287112 510620 287118 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 364334 501004 364340 501016
rect 3292 500976 364340 501004
rect 3292 500964 3298 500976
rect 364334 500964 364340 500976
rect 364392 500964 364398 501016
rect 284294 484372 284300 484424
rect 284352 484412 284358 484424
rect 580166 484412 580172 484424
rect 284352 484384 580172 484412
rect 284352 484372 284358 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 285858 470568 285864 470620
rect 285916 470608 285922 470620
rect 579982 470608 579988 470620
rect 285916 470580 579988 470608
rect 285916 470568 285922 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 104894 468460 104900 468512
rect 104952 468500 104958 468512
rect 339586 468500 339592 468512
rect 104952 468472 339592 468500
rect 104952 468460 104958 468472
rect 339586 468460 339592 468472
rect 339644 468460 339650 468512
rect 169754 467100 169760 467152
rect 169812 467140 169818 467152
rect 334802 467140 334808 467152
rect 169812 467112 334808 467140
rect 169812 467100 169818 467112
rect 334802 467100 334808 467112
rect 334860 467100 334866 467152
rect 299474 465672 299480 465724
rect 299532 465712 299538 465724
rect 325694 465712 325700 465724
rect 299532 465684 325700 465712
rect 299532 465672 299538 465684
rect 325694 465672 325700 465684
rect 325752 465672 325758 465724
rect 316034 464312 316040 464364
rect 316092 464352 316098 464364
rect 429194 464352 429200 464364
rect 316092 464324 429200 464352
rect 316092 464312 316098 464324
rect 429194 464312 429200 464324
rect 429252 464312 429258 464364
rect 226978 462476 226984 462528
rect 227036 462516 227042 462528
rect 375926 462516 375932 462528
rect 227036 462488 375932 462516
rect 227036 462476 227042 462488
rect 375926 462476 375932 462488
rect 375984 462476 375990 462528
rect 225598 462408 225604 462460
rect 225656 462448 225662 462460
rect 380894 462448 380900 462460
rect 225656 462420 380900 462448
rect 225656 462408 225662 462420
rect 380894 462408 380900 462420
rect 380952 462408 380958 462460
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 371234 462380 371240 462392
rect 3568 462352 371240 462380
rect 3568 462340 3574 462352
rect 371234 462340 371240 462352
rect 371292 462340 371298 462392
rect 311802 461592 311808 461644
rect 311860 461632 311866 461644
rect 494054 461632 494060 461644
rect 311860 461604 494060 461632
rect 311860 461592 311866 461604
rect 494054 461592 494060 461604
rect 494112 461592 494118 461644
rect 233970 461320 233976 461372
rect 234028 461360 234034 461372
rect 369854 461360 369860 461372
rect 234028 461332 369860 461360
rect 234028 461320 234034 461332
rect 369854 461320 369860 461332
rect 369912 461320 369918 461372
rect 280062 461252 280068 461304
rect 280120 461292 280126 461304
rect 417510 461292 417516 461304
rect 280120 461264 417516 461292
rect 280120 461252 280126 461264
rect 417510 461252 417516 461264
rect 417568 461252 417574 461304
rect 278682 461184 278688 461236
rect 278740 461224 278746 461236
rect 422938 461224 422944 461236
rect 278740 461196 422944 461224
rect 278740 461184 278746 461196
rect 422938 461184 422944 461196
rect 422996 461184 423002 461236
rect 273990 461116 273996 461168
rect 274048 461156 274054 461168
rect 420178 461156 420184 461168
rect 274048 461128 420184 461156
rect 274048 461116 274054 461128
rect 420178 461116 420184 461128
rect 420236 461116 420242 461168
rect 228358 461048 228364 461100
rect 228416 461088 228422 461100
rect 379146 461088 379152 461100
rect 228416 461060 379152 461088
rect 228416 461048 228422 461060
rect 379146 461048 379152 461060
rect 379204 461048 379210 461100
rect 229738 460980 229744 461032
rect 229796 461020 229802 461032
rect 396534 461020 396540 461032
rect 229796 460992 396540 461020
rect 229796 460980 229802 460992
rect 396534 460980 396540 460992
rect 396592 460980 396598 461032
rect 4890 460912 4896 460964
rect 4948 460952 4954 460964
rect 391934 460952 391940 460964
rect 4948 460924 391940 460952
rect 4948 460912 4954 460924
rect 391934 460912 391940 460924
rect 391992 460912 391998 460964
rect 318150 460844 318156 460896
rect 318208 460884 318214 460896
rect 397454 460884 397460 460896
rect 318208 460856 397460 460884
rect 318208 460844 318214 460856
rect 397454 460844 397460 460856
rect 397512 460844 397518 460896
rect 201494 460776 201500 460828
rect 201552 460816 201558 460828
rect 331766 460816 331772 460828
rect 201552 460788 331772 460816
rect 201552 460776 201558 460788
rect 331766 460776 331772 460788
rect 331824 460776 331830 460828
rect 313090 460708 313096 460760
rect 313148 460748 313154 460760
rect 462314 460748 462320 460760
rect 313148 460720 462320 460748
rect 313148 460708 313154 460720
rect 462314 460708 462320 460720
rect 462372 460708 462378 460760
rect 315022 460640 315028 460692
rect 315080 460680 315086 460692
rect 477494 460680 477500 460692
rect 315080 460652 477500 460680
rect 315080 460640 315086 460652
rect 477494 460640 477500 460652
rect 477552 460640 477558 460692
rect 136634 460572 136640 460624
rect 136692 460612 136698 460624
rect 336734 460612 336740 460624
rect 136692 460584 336740 460612
rect 136692 460572 136698 460584
rect 336734 460572 336740 460584
rect 336792 460572 336798 460624
rect 308674 460504 308680 460556
rect 308732 460544 308738 460556
rect 527174 460544 527180 460556
rect 308732 460516 527180 460544
rect 308732 460504 308738 460516
rect 527174 460504 527180 460516
rect 527232 460504 527238 460556
rect 310238 460436 310244 460488
rect 310296 460476 310302 460488
rect 542354 460476 542360 460488
rect 310296 460448 542360 460476
rect 310296 460436 310302 460448
rect 542354 460436 542360 460448
rect 542412 460436 542418 460488
rect 3602 460368 3608 460420
rect 3660 460408 3666 460420
rect 353846 460408 353852 460420
rect 3660 460380 353852 460408
rect 3660 460368 3666 460380
rect 353846 460368 353852 460380
rect 353904 460368 353910 460420
rect 3694 460300 3700 460352
rect 3752 460340 3758 460352
rect 358814 460340 358820 460352
rect 3752 460312 358820 460340
rect 3752 460300 3758 460312
rect 358814 460300 358820 460312
rect 358872 460300 358878 460352
rect 3786 460232 3792 460284
rect 3844 460272 3850 460284
rect 363322 460272 363328 460284
rect 3844 460244 363328 460272
rect 3844 460232 3850 460244
rect 363322 460232 363328 460244
rect 363380 460232 363386 460284
rect 3878 460164 3884 460216
rect 3936 460204 3942 460216
rect 368106 460204 368112 460216
rect 3936 460176 368112 460204
rect 3936 460164 3942 460176
rect 368106 460164 368112 460176
rect 368164 460164 368170 460216
rect 266354 460096 266360 460148
rect 266412 460136 266418 460148
rect 327074 460136 327080 460148
rect 266412 460108 327080 460136
rect 266412 460096 266418 460108
rect 327074 460096 327080 460108
rect 327132 460096 327138 460148
rect 324130 460028 324136 460080
rect 324188 460068 324194 460080
rect 347774 460068 347780 460080
rect 324188 460040 347780 460068
rect 324188 460028 324194 460040
rect 347774 460028 347780 460040
rect 347832 460028 347838 460080
rect 322842 459960 322848 460012
rect 322900 460000 322906 460012
rect 331214 460000 331220 460012
rect 322900 459972 331220 460000
rect 322900 459960 322906 459972
rect 331214 459960 331220 459972
rect 331272 459960 331278 460012
rect 355962 459552 355968 459604
rect 356020 459592 356026 459604
rect 374362 459592 374368 459604
rect 356020 459564 374368 459592
rect 356020 459552 356026 459564
rect 374362 459552 374368 459564
rect 374420 459552 374426 459604
rect 233878 458804 233884 458856
rect 233936 458844 233942 458856
rect 377582 458844 377588 458856
rect 233936 458816 377588 458844
rect 233936 458804 233942 458816
rect 377582 458804 377588 458816
rect 377640 458804 377646 458856
rect 275554 458736 275560 458788
rect 275612 458776 275618 458788
rect 424318 458776 424324 458788
rect 275612 458748 424324 458776
rect 275612 458736 275618 458748
rect 424318 458736 424324 458748
rect 424376 458736 424382 458788
rect 277118 458668 277124 458720
rect 277176 458708 277182 458720
rect 425698 458708 425704 458720
rect 277176 458680 425704 458708
rect 277176 458668 277182 458680
rect 425698 458668 425704 458680
rect 425756 458668 425762 458720
rect 232498 458600 232504 458652
rect 232556 458640 232562 458652
rect 382274 458640 382280 458652
rect 232556 458612 382280 458640
rect 232556 458600 232562 458612
rect 382274 458600 382280 458612
rect 382332 458600 382338 458652
rect 231118 458532 231124 458584
rect 231176 458572 231182 458584
rect 387058 458572 387064 458584
rect 231176 458544 387064 458572
rect 231176 458532 231182 458544
rect 387058 458532 387064 458544
rect 387116 458532 387122 458584
rect 255038 458464 255044 458516
rect 255096 458504 255102 458516
rect 421558 458504 421564 458516
rect 255096 458476 421564 458504
rect 255096 458464 255102 458476
rect 421558 458464 421564 458476
rect 421616 458464 421622 458516
rect 245562 458396 245568 458448
rect 245620 458436 245626 458448
rect 418798 458436 418804 458448
rect 245620 458408 418804 458436
rect 245620 458396 245626 458408
rect 418798 458396 418804 458408
rect 418856 458396 418862 458448
rect 240778 458328 240784 458380
rect 240836 458368 240842 458380
rect 417418 458368 417424 458380
rect 240836 458340 417424 458368
rect 240836 458328 240842 458340
rect 417418 458328 417424 458340
rect 417476 458328 417482 458380
rect 235902 458260 235908 458312
rect 235960 458300 235966 458312
rect 580258 458300 580264 458312
rect 235960 458272 580264 458300
rect 235960 458260 235966 458272
rect 580258 458260 580264 458272
rect 580316 458260 580322 458312
rect 3510 458192 3516 458244
rect 3568 458232 3574 458244
rect 373120 458232 373126 458244
rect 3568 458204 373126 458232
rect 3568 458192 3574 458204
rect 373120 458192 373126 458204
rect 373178 458192 373184 458244
rect 273226 457660 292574 457688
rect 3418 457444 3424 457496
rect 3476 457484 3482 457496
rect 273226 457484 273254 457660
rect 281626 457580 281632 457632
rect 281684 457620 281690 457632
rect 281684 457592 287836 457620
rect 281684 457580 281690 457592
rect 3476 457456 273254 457484
rect 3476 457444 3482 457456
rect 283374 457444 283380 457496
rect 283432 457444 283438 457496
rect 283392 456804 283420 457444
rect 287808 457416 287836 457592
rect 292546 457484 292574 457660
rect 355962 457484 355968 457496
rect 292546 457456 355968 457484
rect 355962 457444 355968 457456
rect 356020 457444 356026 457496
rect 287808 457388 296714 457416
rect 296686 456872 296714 457388
rect 427078 456872 427084 456884
rect 296686 456844 427084 456872
rect 427078 456832 427084 456844
rect 427136 456832 427142 456884
rect 580166 456804 580172 456816
rect 283392 456776 580172 456804
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 233970 449868 233976 449880
rect 3384 449840 233976 449868
rect 3384 449828 3390 449840
rect 233970 449828 233976 449840
rect 234028 449828 234034 449880
rect 417510 431876 417516 431928
rect 417568 431916 417574 431928
rect 580166 431916 580172 431928
rect 417568 431888 580172 431916
rect 417568 431876 417574 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 427078 419432 427084 419484
rect 427136 419472 427142 419484
rect 580166 419472 580172 419484
rect 427136 419444 580172 419472
rect 427136 419432 427142 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 226978 411244 226984 411256
rect 3016 411216 226984 411244
rect 3016 411204 3022 411216
rect 226978 411204 226984 411216
rect 227036 411204 227042 411256
rect 422938 405628 422944 405680
rect 422996 405668 423002 405680
rect 579614 405668 579620 405680
rect 422996 405640 579620 405668
rect 422996 405628 423002 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 424318 379448 424324 379500
rect 424376 379488 424382 379500
rect 580166 379488 580172 379500
rect 424376 379460 580172 379488
rect 424376 379448 424382 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 233878 372552 233884 372564
rect 3292 372524 233884 372552
rect 3292 372512 3298 372524
rect 233878 372512 233884 372524
rect 233936 372512 233942 372564
rect 425698 365644 425704 365696
rect 425756 365684 425762 365696
rect 580166 365684 580172 365696
rect 425756 365656 580172 365684
rect 425756 365644 425762 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 225598 358748 225604 358760
rect 3384 358720 225604 358748
rect 3384 358708 3390 358720
rect 225598 358708 225604 358720
rect 225656 358708 225662 358760
rect 420178 353200 420184 353252
rect 420236 353240 420242 353252
rect 580166 353240 580172 353252
rect 420236 353212 580172 353240
rect 420236 353200 420242 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 228358 346372 228364 346384
rect 3200 346344 228364 346372
rect 3200 346332 3206 346344
rect 228358 346332 228364 346344
rect 228416 346332 228422 346384
rect 294414 336744 294420 336796
rect 294472 336744 294478 336796
rect 233970 336676 233976 336728
rect 234028 336716 234034 336728
rect 237006 336716 237012 336728
rect 234028 336688 237012 336716
rect 234028 336676 234034 336688
rect 237006 336676 237012 336688
rect 237064 336676 237070 336728
rect 239398 336676 239404 336728
rect 239456 336716 239462 336728
rect 240134 336716 240140 336728
rect 239456 336688 240140 336716
rect 239456 336676 239462 336688
rect 240134 336676 240140 336688
rect 240192 336676 240198 336728
rect 260834 336676 260840 336728
rect 260892 336716 260898 336728
rect 261110 336716 261116 336728
rect 260892 336688 261116 336716
rect 260892 336676 260898 336688
rect 261110 336676 261116 336688
rect 261168 336676 261174 336728
rect 271138 336676 271144 336728
rect 271196 336716 271202 336728
rect 272426 336716 272432 336728
rect 271196 336688 272432 336716
rect 271196 336676 271202 336688
rect 272426 336676 272432 336688
rect 272484 336676 272490 336728
rect 293218 336676 293224 336728
rect 293276 336716 293282 336728
rect 294432 336716 294460 336744
rect 293276 336688 294460 336716
rect 293276 336676 293282 336688
rect 296806 336676 296812 336728
rect 296864 336716 296870 336728
rect 297266 336716 297272 336728
rect 296864 336688 297272 336716
rect 296864 336676 296870 336688
rect 297266 336676 297272 336688
rect 297324 336676 297330 336728
rect 300762 336676 300768 336728
rect 300820 336716 300826 336728
rect 304074 336716 304080 336728
rect 300820 336688 304080 336716
rect 300820 336676 300826 336688
rect 304074 336676 304080 336688
rect 304132 336676 304138 336728
rect 309318 336676 309324 336728
rect 309376 336716 309382 336728
rect 309502 336716 309508 336728
rect 309376 336688 309508 336716
rect 309376 336676 309382 336688
rect 309502 336676 309508 336688
rect 309560 336676 309566 336728
rect 335446 336676 335452 336728
rect 335504 336716 335510 336728
rect 335630 336716 335636 336728
rect 335504 336688 335636 336716
rect 335504 336676 335510 336688
rect 335630 336676 335636 336688
rect 335688 336676 335694 336728
rect 346394 336676 346400 336728
rect 346452 336716 346458 336728
rect 346670 336716 346676 336728
rect 346452 336688 346676 336716
rect 346452 336676 346458 336688
rect 346670 336676 346676 336688
rect 346728 336676 346734 336728
rect 367094 336676 367100 336728
rect 367152 336716 367158 336728
rect 367462 336716 367468 336728
rect 367152 336688 367468 336716
rect 367152 336676 367158 336688
rect 367462 336676 367468 336688
rect 367520 336676 367526 336728
rect 376754 336676 376760 336728
rect 376812 336716 376818 336728
rect 377030 336716 377036 336728
rect 376812 336688 377036 336716
rect 376812 336676 376818 336688
rect 377030 336676 377036 336688
rect 377088 336676 377094 336728
rect 386414 336676 386420 336728
rect 386472 336716 386478 336728
rect 386782 336716 386788 336728
rect 386472 336688 386788 336716
rect 386472 336676 386478 336688
rect 386782 336676 386788 336688
rect 386840 336676 386846 336728
rect 397546 336676 397552 336728
rect 397604 336716 397610 336728
rect 397822 336716 397828 336728
rect 397604 336688 397828 336716
rect 397604 336676 397610 336688
rect 397822 336676 397828 336688
rect 397880 336676 397886 336728
rect 401594 336676 401600 336728
rect 401652 336716 401658 336728
rect 401870 336716 401876 336728
rect 401652 336688 401876 336716
rect 401652 336676 401658 336688
rect 401870 336676 401876 336688
rect 401928 336676 401934 336728
rect 367186 336608 367192 336660
rect 367244 336648 367250 336660
rect 367738 336648 367744 336660
rect 367244 336620 367744 336648
rect 367244 336608 367250 336620
rect 367738 336608 367744 336620
rect 367796 336608 367802 336660
rect 253198 336540 253204 336592
rect 253256 336580 253262 336592
rect 253934 336580 253940 336592
rect 253256 336552 253940 336580
rect 253256 336540 253262 336552
rect 253934 336540 253940 336552
rect 253992 336540 253998 336592
rect 289170 336540 289176 336592
rect 289228 336580 289234 336592
rect 289998 336580 290004 336592
rect 289228 336552 290004 336580
rect 289228 336540 289234 336552
rect 289998 336540 290004 336552
rect 290056 336540 290062 336592
rect 298738 336540 298744 336592
rect 298796 336580 298802 336592
rect 302418 336580 302424 336592
rect 298796 336552 302424 336580
rect 298796 336540 298802 336552
rect 302418 336540 302424 336552
rect 302476 336540 302482 336592
rect 340782 336540 340788 336592
rect 340840 336580 340846 336592
rect 341334 336580 341340 336592
rect 340840 336552 341340 336580
rect 340840 336540 340846 336552
rect 341334 336540 341340 336552
rect 341392 336540 341398 336592
rect 399754 336540 399760 336592
rect 399812 336580 399818 336592
rect 400858 336580 400864 336592
rect 399812 336552 400864 336580
rect 399812 336540 399818 336552
rect 400858 336540 400864 336552
rect 400916 336540 400922 336592
rect 269758 336472 269764 336524
rect 269816 336512 269822 336524
rect 271874 336512 271880 336524
rect 269816 336484 271880 336512
rect 269816 336472 269822 336484
rect 271874 336472 271880 336484
rect 271932 336472 271938 336524
rect 294598 336472 294604 336524
rect 294656 336512 294662 336524
rect 298554 336512 298560 336524
rect 294656 336484 298560 336512
rect 294656 336472 294662 336484
rect 298554 336472 298560 336484
rect 298612 336472 298618 336524
rect 303062 336472 303068 336524
rect 303120 336512 303126 336524
rect 305362 336512 305368 336524
rect 303120 336484 305368 336512
rect 303120 336472 303126 336484
rect 305362 336472 305368 336484
rect 305420 336472 305426 336524
rect 350074 336472 350080 336524
rect 350132 336512 350138 336524
rect 358078 336512 358084 336524
rect 350132 336484 358084 336512
rect 350132 336472 350138 336484
rect 358078 336472 358084 336484
rect 358136 336472 358142 336524
rect 362862 336472 362868 336524
rect 362920 336512 362926 336524
rect 373350 336512 373356 336524
rect 362920 336484 373356 336512
rect 362920 336472 362926 336484
rect 373350 336472 373356 336484
rect 373408 336472 373414 336524
rect 233878 336404 233884 336456
rect 233936 336444 233942 336456
rect 233936 336416 296714 336444
rect 233936 336404 233942 336416
rect 124214 336336 124220 336388
rect 124272 336376 124278 336388
rect 273254 336376 273260 336388
rect 124272 336348 273260 336376
rect 124272 336336 124278 336348
rect 273254 336336 273260 336348
rect 273312 336336 273318 336388
rect 296686 336376 296714 336416
rect 297450 336404 297456 336456
rect 297508 336444 297514 336456
rect 299842 336444 299848 336456
rect 297508 336416 299848 336444
rect 297508 336404 297514 336416
rect 299842 336404 299848 336416
rect 299900 336404 299906 336456
rect 302878 336404 302884 336456
rect 302936 336444 302942 336456
rect 309686 336444 309692 336456
rect 302936 336416 309692 336444
rect 302936 336404 302942 336416
rect 309686 336404 309692 336416
rect 309744 336404 309750 336456
rect 353754 336404 353760 336456
rect 353812 336444 353818 336456
rect 382918 336444 382924 336456
rect 353812 336416 382924 336444
rect 353812 336404 353818 336416
rect 382918 336404 382924 336416
rect 382976 336404 382982 336456
rect 302234 336376 302240 336388
rect 296686 336348 302240 336376
rect 302234 336336 302240 336348
rect 302292 336336 302298 336388
rect 305822 336336 305828 336388
rect 305880 336376 305886 336388
rect 313366 336376 313372 336388
rect 305880 336348 313372 336376
rect 305880 336336 305886 336348
rect 313366 336336 313372 336348
rect 313424 336336 313430 336388
rect 358170 336336 358176 336388
rect 358228 336376 358234 336388
rect 387058 336376 387064 336388
rect 358228 336348 387064 336376
rect 358228 336336 358234 336348
rect 387058 336336 387064 336348
rect 387116 336336 387122 336388
rect 396442 336336 396448 336388
rect 396500 336376 396506 336388
rect 422938 336376 422944 336388
rect 396500 336348 422944 336376
rect 396500 336336 396506 336348
rect 422938 336336 422944 336348
rect 422996 336336 423002 336388
rect 117314 336268 117320 336320
rect 117372 336308 117378 336320
rect 271046 336308 271052 336320
rect 117372 336280 271052 336308
rect 117372 336268 117378 336280
rect 271046 336268 271052 336280
rect 271104 336268 271110 336320
rect 286410 336268 286416 336320
rect 286468 336308 286474 336320
rect 287790 336308 287796 336320
rect 286468 336280 287796 336308
rect 286468 336268 286474 336280
rect 287790 336268 287796 336280
rect 287848 336268 287854 336320
rect 302970 336268 302976 336320
rect 303028 336308 303034 336320
rect 314838 336308 314844 336320
rect 303028 336280 314844 336308
rect 303028 336268 303034 336280
rect 314838 336268 314844 336280
rect 314896 336268 314902 336320
rect 315298 336268 315304 336320
rect 315356 336308 315362 336320
rect 324314 336308 324320 336320
rect 315356 336280 324320 336308
rect 315356 336268 315362 336280
rect 324314 336268 324320 336280
rect 324372 336268 324378 336320
rect 334342 336268 334348 336320
rect 334400 336308 334406 336320
rect 338206 336308 338212 336320
rect 334400 336280 338212 336308
rect 334400 336268 334406 336280
rect 338206 336268 338212 336280
rect 338264 336268 338270 336320
rect 343818 336268 343824 336320
rect 343876 336308 343882 336320
rect 345658 336308 345664 336320
rect 343876 336280 345664 336308
rect 343876 336268 343882 336280
rect 345658 336268 345664 336280
rect 345716 336268 345722 336320
rect 345750 336268 345756 336320
rect 345808 336308 345814 336320
rect 357434 336308 357440 336320
rect 345808 336280 357440 336308
rect 345808 336268 345814 336280
rect 357434 336268 357440 336280
rect 357492 336268 357498 336320
rect 362770 336268 362776 336320
rect 362828 336308 362834 336320
rect 370498 336308 370504 336320
rect 362828 336280 370504 336308
rect 362828 336268 362834 336280
rect 370498 336268 370504 336280
rect 370556 336268 370562 336320
rect 373074 336268 373080 336320
rect 373132 336308 373138 336320
rect 447134 336308 447140 336320
rect 373132 336280 447140 336308
rect 373132 336268 373138 336280
rect 447134 336268 447140 336280
rect 447192 336268 447198 336320
rect 110414 336200 110420 336252
rect 110472 336240 110478 336252
rect 268838 336240 268844 336252
rect 110472 336212 268844 336240
rect 110472 336200 110478 336212
rect 268838 336200 268844 336212
rect 268896 336200 268902 336252
rect 307018 336200 307024 336252
rect 307076 336240 307082 336252
rect 322106 336240 322112 336252
rect 307076 336212 322112 336240
rect 307076 336200 307082 336212
rect 322106 336200 322112 336212
rect 322164 336200 322170 336252
rect 339494 336200 339500 336252
rect 339552 336240 339558 336252
rect 339678 336240 339684 336252
rect 339552 336212 339684 336240
rect 339552 336200 339558 336212
rect 339678 336200 339684 336212
rect 339736 336200 339742 336252
rect 347314 336200 347320 336252
rect 347372 336240 347378 336252
rect 362954 336240 362960 336252
rect 347372 336212 362960 336240
rect 347372 336200 347378 336212
rect 362954 336200 362960 336212
rect 363012 336200 363018 336252
rect 375282 336200 375288 336252
rect 375340 336240 375346 336252
rect 454034 336240 454040 336252
rect 375340 336212 454040 336240
rect 375340 336200 375346 336212
rect 454034 336200 454040 336212
rect 454092 336200 454098 336252
rect 99374 336132 99380 336184
rect 99432 336172 99438 336184
rect 265526 336172 265532 336184
rect 99432 336144 265532 336172
rect 99432 336132 99438 336144
rect 265526 336132 265532 336144
rect 265584 336132 265590 336184
rect 297358 336132 297364 336184
rect 297416 336172 297422 336184
rect 311894 336172 311900 336184
rect 297416 336144 311900 336172
rect 297416 336132 297422 336144
rect 311894 336132 311900 336144
rect 311952 336132 311958 336184
rect 324314 336132 324320 336184
rect 324372 336172 324378 336184
rect 334894 336172 334900 336184
rect 324372 336144 334900 336172
rect 324372 336132 324378 336144
rect 334894 336132 334900 336144
rect 334952 336132 334958 336184
rect 348602 336132 348608 336184
rect 348660 336172 348666 336184
rect 359458 336172 359464 336184
rect 348660 336144 359464 336172
rect 348660 336132 348666 336144
rect 359458 336132 359464 336144
rect 359516 336132 359522 336184
rect 377490 336132 377496 336184
rect 377548 336172 377554 336184
rect 460934 336172 460940 336184
rect 377548 336144 460940 336172
rect 377548 336132 377554 336144
rect 460934 336132 460940 336144
rect 460992 336132 460998 336184
rect 15838 336064 15844 336116
rect 15896 336104 15902 336116
rect 238110 336104 238116 336116
rect 15896 336076 238116 336104
rect 15896 336064 15902 336076
rect 238110 336064 238116 336076
rect 238168 336064 238174 336116
rect 276658 336064 276664 336116
rect 276716 336104 276722 336116
rect 285674 336104 285680 336116
rect 276716 336076 285680 336104
rect 276716 336064 276722 336076
rect 285674 336064 285680 336076
rect 285732 336064 285738 336116
rect 289078 336064 289084 336116
rect 289136 336104 289142 336116
rect 310790 336104 310796 336116
rect 289136 336076 310796 336104
rect 289136 336064 289142 336076
rect 310790 336064 310796 336076
rect 310848 336064 310854 336116
rect 327074 336064 327080 336116
rect 327132 336104 327138 336116
rect 335998 336104 336004 336116
rect 327132 336076 336004 336104
rect 327132 336064 327138 336076
rect 335998 336064 336004 336076
rect 336056 336064 336062 336116
rect 350810 336064 350816 336116
rect 350868 336104 350874 336116
rect 373994 336104 374000 336116
rect 350868 336076 374000 336104
rect 350868 336064 350874 336076
rect 373994 336064 374000 336076
rect 374052 336064 374058 336116
rect 379882 336064 379888 336116
rect 379940 336104 379946 336116
rect 467834 336104 467840 336116
rect 379940 336076 467840 336104
rect 379940 336064 379946 336076
rect 467834 336064 467840 336076
rect 467892 336064 467898 336116
rect 6178 335996 6184 336048
rect 6236 336036 6242 336048
rect 236270 336036 236276 336048
rect 6236 336008 236276 336036
rect 6236 335996 6242 336008
rect 236270 335996 236276 336008
rect 236328 335996 236334 336048
rect 269298 335996 269304 336048
rect 269356 336036 269362 336048
rect 284478 336036 284484 336048
rect 269356 336008 284484 336036
rect 269356 335996 269362 336008
rect 284478 335996 284484 336008
rect 284536 335996 284542 336048
rect 286226 335996 286232 336048
rect 286284 336036 286290 336048
rect 291194 336036 291200 336048
rect 286284 336008 291200 336036
rect 286284 335996 286290 336008
rect 291194 335996 291200 336008
rect 291252 335996 291258 336048
rect 315206 336036 315212 336048
rect 296686 336008 315212 336036
rect 264238 335928 264244 335980
rect 264296 335968 264302 335980
rect 266998 335968 267004 335980
rect 264296 335940 267004 335968
rect 264296 335928 264302 335940
rect 266998 335928 267004 335940
rect 267056 335928 267062 335980
rect 291838 335928 291844 335980
rect 291896 335968 291902 335980
rect 296686 335968 296714 336008
rect 315206 335996 315212 336008
rect 315264 335996 315270 336048
rect 320174 335996 320180 336048
rect 320232 336036 320238 336048
rect 333974 336036 333980 336048
rect 320232 336008 333980 336036
rect 320232 335996 320238 336008
rect 333974 335996 333980 336008
rect 334032 335996 334038 336048
rect 344922 335996 344928 336048
rect 344980 336036 344986 336048
rect 351178 336036 351184 336048
rect 344980 336008 351184 336036
rect 344980 335996 344986 336008
rect 351178 335996 351184 336008
rect 351236 335996 351242 336048
rect 351914 335996 351920 336048
rect 351972 336036 351978 336048
rect 377398 336036 377404 336048
rect 351972 336008 377404 336036
rect 351972 335996 351978 336008
rect 377398 335996 377404 336008
rect 377456 335996 377462 336048
rect 381814 335996 381820 336048
rect 381872 336036 381878 336048
rect 474734 336036 474740 336048
rect 381872 336008 474740 336036
rect 381872 335996 381878 336008
rect 474734 335996 474740 336008
rect 474792 335996 474798 336048
rect 291896 335940 296714 335968
rect 291896 335928 291902 335940
rect 305638 335928 305644 335980
rect 305696 335968 305702 335980
rect 307202 335968 307208 335980
rect 305696 335940 307208 335968
rect 305696 335928 305702 335940
rect 307202 335928 307208 335940
rect 307260 335928 307266 335980
rect 359458 335928 359464 335980
rect 359516 335968 359522 335980
rect 366174 335968 366180 335980
rect 359516 335940 366180 335968
rect 359516 335928 359522 335940
rect 366174 335928 366180 335940
rect 366232 335928 366238 335980
rect 251818 335860 251824 335912
rect 251876 335900 251882 335912
rect 253014 335900 253020 335912
rect 251876 335872 253020 335900
rect 251876 335860 251882 335872
rect 253014 335860 253020 335872
rect 253072 335860 253078 335912
rect 291930 335792 291936 335844
rect 291988 335832 291994 335844
rect 293310 335832 293316 335844
rect 291988 335804 293316 335832
rect 291988 335792 291994 335804
rect 293310 335792 293316 335804
rect 293368 335792 293374 335844
rect 319438 335792 319444 335844
rect 319496 335832 319502 335844
rect 321002 335832 321008 335844
rect 319496 335804 321008 335832
rect 319496 335792 319502 335804
rect 321002 335792 321008 335804
rect 321060 335792 321066 335844
rect 273898 335724 273904 335776
rect 273956 335764 273962 335776
rect 277946 335764 277952 335776
rect 273956 335736 277952 335764
rect 273956 335724 273962 335736
rect 277946 335724 277952 335736
rect 278004 335724 278010 335776
rect 287698 335656 287704 335708
rect 287756 335696 287762 335708
rect 290366 335696 290372 335708
rect 287756 335668 290372 335696
rect 287756 335656 287762 335668
rect 290366 335656 290372 335668
rect 290424 335656 290430 335708
rect 322198 335656 322204 335708
rect 322256 335696 322262 335708
rect 326522 335696 326528 335708
rect 322256 335668 326528 335696
rect 322256 335656 322262 335668
rect 326522 335656 326528 335668
rect 326580 335656 326586 335708
rect 340966 335656 340972 335708
rect 341024 335696 341030 335708
rect 342254 335696 342260 335708
rect 341024 335668 342260 335696
rect 341024 335656 341030 335668
rect 342254 335656 342260 335668
rect 342312 335656 342318 335708
rect 244918 335520 244924 335572
rect 244976 335560 244982 335572
rect 246206 335560 246212 335572
rect 244976 335532 246212 335560
rect 244976 335520 244982 335532
rect 246206 335520 246212 335532
rect 246264 335520 246270 335572
rect 301498 335452 301504 335504
rect 301556 335492 301562 335504
rect 308582 335492 308588 335504
rect 301556 335464 308588 335492
rect 301556 335452 301562 335464
rect 308582 335452 308588 335464
rect 308640 335452 308646 335504
rect 320818 335452 320824 335504
rect 320876 335492 320882 335504
rect 327626 335492 327632 335504
rect 320876 335464 327632 335492
rect 320876 335452 320882 335464
rect 327626 335452 327632 335464
rect 327684 335452 327690 335504
rect 361758 335452 361764 335504
rect 361816 335492 361822 335504
rect 364978 335492 364984 335504
rect 361816 335464 364984 335492
rect 361816 335452 361822 335464
rect 364978 335452 364984 335464
rect 365036 335452 365042 335504
rect 379974 335384 379980 335436
rect 380032 335424 380038 335436
rect 381538 335424 381544 335436
rect 380032 335396 381544 335424
rect 380032 335384 380038 335396
rect 381538 335384 381544 335396
rect 381596 335384 381602 335436
rect 295978 335316 295984 335368
rect 296036 335356 296042 335368
rect 296714 335356 296720 335368
rect 296036 335328 296720 335356
rect 296036 335316 296042 335328
rect 296714 335316 296720 335328
rect 296772 335316 296778 335368
rect 304258 335316 304264 335368
rect 304316 335356 304322 335368
rect 307846 335356 307852 335368
rect 304316 335328 307852 335356
rect 304316 335316 304322 335328
rect 307846 335316 307852 335328
rect 307904 335316 307910 335368
rect 313918 335316 313924 335368
rect 313976 335356 313982 335368
rect 317414 335356 317420 335368
rect 313976 335328 317420 335356
rect 313976 335316 313982 335328
rect 317414 335316 317420 335328
rect 317472 335316 317478 335368
rect 333238 335316 333244 335368
rect 333296 335356 333302 335368
rect 337102 335356 337108 335368
rect 333296 335328 337108 335356
rect 333296 335316 333302 335328
rect 337102 335316 337108 335328
rect 337160 335316 337166 335368
rect 402330 335316 402336 335368
rect 402388 335356 402394 335368
rect 403618 335356 403624 335368
rect 402388 335328 403624 335356
rect 402388 335316 402394 335328
rect 403618 335316 403624 335328
rect 403676 335316 403682 335368
rect 411806 335316 411812 335368
rect 411864 335356 411870 335368
rect 413370 335356 413376 335368
rect 411864 335328 413376 335356
rect 411864 335316 411870 335328
rect 413370 335316 413376 335328
rect 413428 335316 413434 335368
rect 321646 335180 321652 335232
rect 321704 335220 321710 335232
rect 321830 335220 321836 335232
rect 321704 335192 321836 335220
rect 321704 335180 321710 335192
rect 321830 335180 321836 335192
rect 321888 335180 321894 335232
rect 383562 334636 383568 334688
rect 383620 334676 383626 334688
rect 480254 334676 480260 334688
rect 383620 334648 480260 334676
rect 383620 334636 383626 334648
rect 480254 334636 480260 334648
rect 480312 334636 480318 334688
rect 224954 334568 224960 334620
rect 225012 334608 225018 334620
rect 300762 334608 300768 334620
rect 225012 334580 300768 334608
rect 225012 334568 225018 334580
rect 300762 334568 300768 334580
rect 300820 334568 300826 334620
rect 403158 334568 403164 334620
rect 403216 334608 403222 334620
rect 543734 334608 543740 334620
rect 403216 334580 543740 334608
rect 403216 334568 403222 334580
rect 543734 334568 543740 334580
rect 543792 334568 543798 334620
rect 414014 334500 414020 334552
rect 414072 334540 414078 334552
rect 414198 334540 414204 334552
rect 414072 334512 414204 334540
rect 414072 334500 414078 334512
rect 414198 334500 414204 334512
rect 414256 334500 414262 334552
rect 384482 333276 384488 333328
rect 384540 333316 384546 333328
rect 483014 333316 483020 333328
rect 384540 333288 483020 333316
rect 384540 333276 384546 333288
rect 483014 333276 483020 333288
rect 483072 333276 483078 333328
rect 227714 333208 227720 333260
rect 227772 333248 227778 333260
rect 303062 333248 303068 333260
rect 227772 333220 303068 333248
rect 227772 333208 227778 333220
rect 303062 333208 303068 333220
rect 303120 333208 303126 333260
rect 408494 333208 408500 333260
rect 408552 333248 408558 333260
rect 561674 333248 561680 333260
rect 408552 333220 561680 333248
rect 408552 333208 408558 333220
rect 561674 333208 561680 333220
rect 561732 333208 561738 333260
rect 175274 331916 175280 331968
rect 175332 331956 175338 331968
rect 288894 331956 288900 331968
rect 175332 331928 288900 331956
rect 175332 331916 175338 331928
rect 288894 331916 288900 331928
rect 288952 331916 288958 331968
rect 390002 331916 390008 331968
rect 390060 331956 390066 331968
rect 500954 331956 500960 331968
rect 390060 331928 500960 331956
rect 390060 331916 390066 331928
rect 500954 331916 500960 331928
rect 501012 331916 501018 331968
rect 46934 331848 46940 331900
rect 46992 331888 46998 331900
rect 249426 331888 249432 331900
rect 46992 331860 249432 331888
rect 46992 331848 46998 331860
rect 249426 331848 249432 331860
rect 249484 331848 249490 331900
rect 403802 331848 403808 331900
rect 403860 331888 403866 331900
rect 546494 331888 546500 331900
rect 403860 331860 546500 331888
rect 403860 331848 403866 331860
rect 546494 331848 546500 331860
rect 546552 331848 546558 331900
rect 383838 331168 383844 331220
rect 383896 331208 383902 331220
rect 384022 331208 384028 331220
rect 383896 331180 384028 331208
rect 383896 331168 383902 331180
rect 384022 331168 384028 331180
rect 384080 331168 384086 331220
rect 347958 330760 347964 330812
rect 348016 330760 348022 330812
rect 238754 330624 238760 330676
rect 238812 330664 238818 330676
rect 239582 330664 239588 330676
rect 238812 330636 239588 330664
rect 238812 330624 238818 330636
rect 239582 330624 239588 330636
rect 239640 330624 239646 330676
rect 347976 330608 348004 330760
rect 168374 330556 168380 330608
rect 168432 330596 168438 330608
rect 286686 330596 286692 330608
rect 168432 330568 286692 330596
rect 168432 330556 168438 330568
rect 286686 330556 286692 330568
rect 286744 330556 286750 330608
rect 347958 330556 347964 330608
rect 348016 330556 348022 330608
rect 366266 330556 366272 330608
rect 366324 330596 366330 330608
rect 423674 330596 423680 330608
rect 366324 330568 423680 330596
rect 366324 330556 366330 330568
rect 423674 330556 423680 330568
rect 423732 330556 423738 330608
rect 57974 330488 57980 330540
rect 58032 330528 58038 330540
rect 58032 330500 238754 330528
rect 58032 330488 58038 330500
rect 234614 330420 234620 330472
rect 234672 330460 234678 330472
rect 235534 330460 235540 330472
rect 234672 330432 235540 330460
rect 234672 330420 234678 330432
rect 235534 330420 235540 330432
rect 235592 330420 235598 330472
rect 238726 330392 238754 330500
rect 238846 330488 238852 330540
rect 238904 330528 238910 330540
rect 239214 330528 239220 330540
rect 238904 330500 239220 330528
rect 238904 330488 238910 330500
rect 239214 330488 239220 330500
rect 239272 330488 239278 330540
rect 240226 330488 240232 330540
rect 240284 330528 240290 330540
rect 240686 330528 240692 330540
rect 240284 330500 240692 330528
rect 240284 330488 240290 330500
rect 240686 330488 240692 330500
rect 240744 330488 240750 330540
rect 241514 330488 241520 330540
rect 241572 330528 241578 330540
rect 242158 330528 242164 330540
rect 241572 330500 242164 330528
rect 241572 330488 241578 330500
rect 242158 330488 242164 330500
rect 242216 330488 242222 330540
rect 243078 330488 243084 330540
rect 243136 330528 243142 330540
rect 243998 330528 244004 330540
rect 243136 330500 244004 330528
rect 243136 330488 243142 330500
rect 243998 330488 244004 330500
rect 244056 330488 244062 330540
rect 254118 330488 254124 330540
rect 254176 330528 254182 330540
rect 254946 330528 254952 330540
rect 254176 330500 254952 330528
rect 254176 330488 254182 330500
rect 254946 330488 254952 330500
rect 255004 330488 255010 330540
rect 255406 330488 255412 330540
rect 255464 330528 255470 330540
rect 255682 330528 255688 330540
rect 255464 330500 255688 330528
rect 255464 330488 255470 330500
rect 255682 330488 255688 330500
rect 255740 330488 255746 330540
rect 256694 330488 256700 330540
rect 256752 330528 256758 330540
rect 257154 330528 257160 330540
rect 256752 330500 257160 330528
rect 256752 330488 256758 330500
rect 257154 330488 257160 330500
rect 257212 330488 257218 330540
rect 258166 330488 258172 330540
rect 258224 330528 258230 330540
rect 258626 330528 258632 330540
rect 258224 330500 258632 330528
rect 258224 330488 258230 330500
rect 258626 330488 258632 330500
rect 258684 330488 258690 330540
rect 259454 330488 259460 330540
rect 259512 330528 259518 330540
rect 260374 330528 260380 330540
rect 259512 330500 260380 330528
rect 259512 330488 259518 330500
rect 260374 330488 260380 330500
rect 260432 330488 260438 330540
rect 260926 330488 260932 330540
rect 260984 330528 260990 330540
rect 261846 330528 261852 330540
rect 260984 330500 261852 330528
rect 260984 330488 260990 330500
rect 261846 330488 261852 330500
rect 261904 330488 261910 330540
rect 262214 330488 262220 330540
rect 262272 330528 262278 330540
rect 262950 330528 262956 330540
rect 262272 330500 262956 330528
rect 262272 330488 262278 330500
rect 262950 330488 262956 330500
rect 263008 330488 263014 330540
rect 265066 330488 265072 330540
rect 265124 330528 265130 330540
rect 265894 330528 265900 330540
rect 265124 330500 265900 330528
rect 265124 330488 265130 330500
rect 265894 330488 265900 330500
rect 265952 330488 265958 330540
rect 266446 330488 266452 330540
rect 266504 330528 266510 330540
rect 267366 330528 267372 330540
rect 266504 330500 267372 330528
rect 266504 330488 266510 330500
rect 267366 330488 267372 330500
rect 267424 330488 267430 330540
rect 267826 330488 267832 330540
rect 267884 330528 267890 330540
rect 268286 330528 268292 330540
rect 267884 330500 268292 330528
rect 267884 330488 267890 330500
rect 268286 330488 268292 330500
rect 268344 330488 268350 330540
rect 269114 330488 269120 330540
rect 269172 330528 269178 330540
rect 269942 330528 269948 330540
rect 269172 330500 269948 330528
rect 269172 330488 269178 330500
rect 269942 330488 269948 330500
rect 270000 330488 270006 330540
rect 270770 330488 270776 330540
rect 270828 330528 270834 330540
rect 271322 330528 271328 330540
rect 270828 330500 271328 330528
rect 270828 330488 270834 330500
rect 271322 330488 271328 330500
rect 271380 330488 271386 330540
rect 271966 330488 271972 330540
rect 272024 330528 272030 330540
rect 272794 330528 272800 330540
rect 272024 330500 272800 330528
rect 272024 330488 272030 330500
rect 272794 330488 272800 330500
rect 272852 330488 272858 330540
rect 285766 330488 285772 330540
rect 285824 330528 285830 330540
rect 286318 330528 286324 330540
rect 285824 330500 286324 330528
rect 285824 330488 285830 330500
rect 286318 330488 286324 330500
rect 286376 330488 286382 330540
rect 291378 330488 291384 330540
rect 291436 330528 291442 330540
rect 292206 330528 292212 330540
rect 291436 330500 292212 330528
rect 291436 330488 291442 330500
rect 292206 330488 292212 330500
rect 292264 330488 292270 330540
rect 302326 330488 302332 330540
rect 302384 330528 302390 330540
rect 303154 330528 303160 330540
rect 302384 330500 303160 330528
rect 302384 330488 302390 330500
rect 303154 330488 303160 330500
rect 303212 330488 303218 330540
rect 305086 330488 305092 330540
rect 305144 330528 305150 330540
rect 305730 330528 305736 330540
rect 305144 330500 305736 330528
rect 305144 330488 305150 330500
rect 305730 330488 305736 330500
rect 305788 330488 305794 330540
rect 306650 330488 306656 330540
rect 306708 330528 306714 330540
rect 307478 330528 307484 330540
rect 306708 330500 307484 330528
rect 306708 330488 306714 330500
rect 307478 330488 307484 330500
rect 307536 330488 307542 330540
rect 309226 330488 309232 330540
rect 309284 330528 309290 330540
rect 310054 330528 310060 330540
rect 309284 330500 310060 330528
rect 309284 330488 309290 330500
rect 310054 330488 310060 330500
rect 310112 330488 310118 330540
rect 310606 330488 310612 330540
rect 310664 330528 310670 330540
rect 311158 330528 311164 330540
rect 310664 330500 311164 330528
rect 310664 330488 310670 330500
rect 311158 330488 311164 330500
rect 311216 330488 311222 330540
rect 313366 330488 313372 330540
rect 313424 330528 313430 330540
rect 314102 330528 314108 330540
rect 313424 330500 314108 330528
rect 313424 330488 313430 330500
rect 314102 330488 314108 330500
rect 314160 330488 314166 330540
rect 314838 330488 314844 330540
rect 314896 330528 314902 330540
rect 315574 330528 315580 330540
rect 314896 330500 315580 330528
rect 314896 330488 314902 330500
rect 315574 330488 315580 330500
rect 315632 330488 315638 330540
rect 316218 330488 316224 330540
rect 316276 330528 316282 330540
rect 316678 330528 316684 330540
rect 316276 330500 316684 330528
rect 316276 330488 316282 330500
rect 316678 330488 316684 330500
rect 316736 330488 316742 330540
rect 318794 330488 318800 330540
rect 318852 330528 318858 330540
rect 319254 330528 319260 330540
rect 318852 330500 319260 330528
rect 318852 330488 318858 330500
rect 319254 330488 319260 330500
rect 319312 330488 319318 330540
rect 331214 330488 331220 330540
rect 331272 330528 331278 330540
rect 331950 330528 331956 330540
rect 331272 330500 331956 330528
rect 331272 330488 331278 330500
rect 331950 330488 331956 330500
rect 332008 330488 332014 330540
rect 332594 330488 332600 330540
rect 332652 330528 332658 330540
rect 333422 330528 333428 330540
rect 332652 330500 333428 330528
rect 332652 330488 332658 330500
rect 333422 330488 333428 330500
rect 333480 330488 333486 330540
rect 334066 330488 334072 330540
rect 334124 330528 334130 330540
rect 334526 330528 334532 330540
rect 334124 330500 334532 330528
rect 334124 330488 334130 330500
rect 334526 330488 334532 330500
rect 334584 330488 334590 330540
rect 336826 330488 336832 330540
rect 336884 330528 336890 330540
rect 337838 330528 337844 330540
rect 336884 330500 337844 330528
rect 336884 330488 336890 330500
rect 337838 330488 337844 330500
rect 337896 330488 337902 330540
rect 342530 330488 342536 330540
rect 342588 330528 342594 330540
rect 342990 330528 342996 330540
rect 342588 330500 342996 330528
rect 342588 330488 342594 330500
rect 342990 330488 342996 330500
rect 343048 330488 343054 330540
rect 345014 330488 345020 330540
rect 345072 330528 345078 330540
rect 345842 330528 345848 330540
rect 345072 330500 345848 330528
rect 345072 330488 345078 330500
rect 345842 330488 345848 330500
rect 345900 330488 345906 330540
rect 347866 330488 347872 330540
rect 347924 330528 347930 330540
rect 348786 330528 348792 330540
rect 347924 330500 348792 330528
rect 347924 330488 347930 330500
rect 348786 330488 348792 330500
rect 348844 330488 348850 330540
rect 360194 330488 360200 330540
rect 360252 330528 360258 330540
rect 360838 330528 360844 330540
rect 360252 330500 360844 330528
rect 360252 330488 360258 330500
rect 360838 330488 360844 330500
rect 360896 330488 360902 330540
rect 364426 330488 364432 330540
rect 364484 330528 364490 330540
rect 365254 330528 365260 330540
rect 364484 330500 365260 330528
rect 364484 330488 364490 330500
rect 365254 330488 365260 330500
rect 365312 330488 365318 330540
rect 367278 330488 367284 330540
rect 367336 330528 367342 330540
rect 368106 330528 368112 330540
rect 367336 330500 368112 330528
rect 367336 330488 367342 330500
rect 368106 330488 368112 330500
rect 368164 330488 368170 330540
rect 368566 330488 368572 330540
rect 368624 330528 368630 330540
rect 369578 330528 369584 330540
rect 368624 330500 369584 330528
rect 368624 330488 368630 330500
rect 369578 330488 369584 330500
rect 369636 330488 369642 330540
rect 390738 330488 390744 330540
rect 390796 330528 390802 330540
rect 391198 330528 391204 330540
rect 390796 330500 391204 330528
rect 390796 330488 390802 330500
rect 391198 330488 391204 330500
rect 391256 330488 391262 330540
rect 392026 330488 392032 330540
rect 392084 330528 392090 330540
rect 392578 330528 392584 330540
rect 392084 330500 392584 330528
rect 392084 330488 392090 330500
rect 392578 330488 392584 330500
rect 392636 330488 392642 330540
rect 393406 330488 393412 330540
rect 393464 330528 393470 330540
rect 394418 330528 394424 330540
rect 393464 330500 394424 330528
rect 393464 330488 393470 330500
rect 394418 330488 394424 330500
rect 394476 330488 394482 330540
rect 396074 330488 396080 330540
rect 396132 330528 396138 330540
rect 396626 330528 396632 330540
rect 396132 330500 396632 330528
rect 396132 330488 396138 330500
rect 396626 330488 396632 330500
rect 396684 330488 396690 330540
rect 397638 330488 397644 330540
rect 397696 330528 397702 330540
rect 398466 330528 398472 330540
rect 397696 330500 398472 330528
rect 397696 330488 397702 330500
rect 398466 330488 398472 330500
rect 398524 330488 398530 330540
rect 550634 330528 550640 330540
rect 408466 330500 550640 330528
rect 255314 330420 255320 330472
rect 255372 330460 255378 330472
rect 256418 330460 256424 330472
rect 255372 330432 256424 330460
rect 255372 330420 255378 330432
rect 256418 330420 256424 330432
rect 256476 330420 256482 330472
rect 256786 330420 256792 330472
rect 256844 330460 256850 330472
rect 257522 330460 257528 330472
rect 256844 330432 257528 330460
rect 256844 330420 256850 330432
rect 257522 330420 257528 330432
rect 257580 330420 257586 330472
rect 258258 330420 258264 330472
rect 258316 330460 258322 330472
rect 258994 330460 259000 330472
rect 258316 330432 259000 330460
rect 258316 330420 258322 330432
rect 258994 330420 259000 330432
rect 259052 330420 259058 330472
rect 262306 330420 262312 330472
rect 262364 330460 262370 330472
rect 263318 330460 263324 330472
rect 262364 330432 263324 330460
rect 262364 330420 262370 330432
rect 263318 330420 263324 330432
rect 263376 330420 263382 330472
rect 316034 330420 316040 330472
rect 316092 330460 316098 330472
rect 317046 330460 317052 330472
rect 316092 330432 317052 330460
rect 316092 330420 316098 330432
rect 317046 330420 317052 330432
rect 317104 330420 317110 330472
rect 331306 330420 331312 330472
rect 331364 330460 331370 330472
rect 332318 330460 332324 330472
rect 331364 330432 332324 330460
rect 331364 330420 331370 330432
rect 332318 330420 332324 330432
rect 332376 330420 332382 330472
rect 342438 330420 342444 330472
rect 342496 330460 342502 330472
rect 343266 330460 343272 330472
rect 342496 330432 343272 330460
rect 342496 330420 342502 330432
rect 343266 330420 343272 330432
rect 343324 330420 343330 330472
rect 390554 330420 390560 330472
rect 390612 330460 390618 330472
rect 391474 330460 391480 330472
rect 390612 330432 391480 330460
rect 390612 330420 390618 330432
rect 391474 330420 391480 330432
rect 391532 330420 391538 330472
rect 391934 330420 391940 330472
rect 391992 330460 391998 330472
rect 392946 330460 392952 330472
rect 391992 330432 392952 330460
rect 391992 330420 391998 330432
rect 392946 330420 392952 330432
rect 393004 330420 393010 330472
rect 396166 330420 396172 330472
rect 396224 330460 396230 330472
rect 396994 330460 397000 330472
rect 396224 330432 397000 330460
rect 396224 330420 396230 330432
rect 396994 330420 397000 330432
rect 397052 330420 397058 330472
rect 397454 330420 397460 330472
rect 397512 330460 397518 330472
rect 398098 330460 398104 330472
rect 397512 330432 398104 330460
rect 397512 330420 397518 330432
rect 398098 330420 398104 330432
rect 398156 330420 398162 330472
rect 252738 330392 252744 330404
rect 238726 330364 252744 330392
rect 252738 330352 252744 330364
rect 252796 330352 252802 330404
rect 405274 330352 405280 330404
rect 405332 330392 405338 330404
rect 408466 330392 408494 330500
rect 550634 330488 550640 330500
rect 550692 330488 550698 330540
rect 405332 330364 408494 330392
rect 405332 330352 405338 330364
rect 258074 330284 258080 330336
rect 258132 330324 258138 330336
rect 258442 330324 258448 330336
rect 258132 330296 258448 330324
rect 258132 330284 258138 330296
rect 258442 330284 258448 330296
rect 258500 330284 258506 330336
rect 317506 330284 317512 330336
rect 317564 330324 317570 330336
rect 318518 330324 318524 330336
rect 317564 330296 318524 330324
rect 317564 330284 317570 330296
rect 318518 330284 318524 330296
rect 318576 330284 318582 330336
rect 287146 330080 287152 330132
rect 287204 330120 287210 330132
rect 288158 330120 288164 330132
rect 287204 330092 288164 330120
rect 287204 330080 287210 330092
rect 288158 330080 288164 330092
rect 288216 330080 288222 330132
rect 394694 329876 394700 329928
rect 394752 329916 394758 329928
rect 395154 329916 395160 329928
rect 394752 329888 395160 329916
rect 394752 329876 394758 329888
rect 395154 329876 395160 329888
rect 395212 329876 395218 329928
rect 340966 329808 340972 329860
rect 341024 329848 341030 329860
rect 341886 329848 341892 329860
rect 341024 329820 341892 329848
rect 341024 329808 341030 329820
rect 341886 329808 341892 329820
rect 341944 329808 341950 329860
rect 241606 329672 241612 329724
rect 241664 329712 241670 329724
rect 242526 329712 242532 329724
rect 241664 329684 242532 329712
rect 241664 329672 241670 329684
rect 242526 329672 242532 329684
rect 242584 329672 242590 329724
rect 267918 329672 267924 329724
rect 267976 329712 267982 329724
rect 268470 329712 268476 329724
rect 267976 329684 268476 329712
rect 267976 329672 267982 329684
rect 268470 329672 268476 329684
rect 268528 329672 268534 329724
rect 365806 329536 365812 329588
rect 365864 329576 365870 329588
rect 366726 329576 366732 329588
rect 365864 329548 366732 329576
rect 365864 329536 365870 329548
rect 366726 329536 366732 329548
rect 366784 329536 366790 329588
rect 201494 329196 201500 329248
rect 201552 329236 201558 329248
rect 296898 329236 296904 329248
rect 201552 329208 296904 329236
rect 201552 329196 201558 329208
rect 296898 329196 296904 329208
rect 296956 329196 296962 329248
rect 160094 329128 160100 329180
rect 160152 329168 160158 329180
rect 269298 329168 269304 329180
rect 160152 329140 269304 329168
rect 160152 329128 160158 329140
rect 269298 329128 269304 329140
rect 269356 329128 269362 329180
rect 26234 329060 26240 329112
rect 26292 329100 26298 329112
rect 242894 329100 242900 329112
rect 26292 329072 242900 329100
rect 26292 329060 26298 329072
rect 242894 329060 242900 329072
rect 242952 329060 242958 329112
rect 392118 329060 392124 329112
rect 392176 329100 392182 329112
rect 507854 329100 507860 329112
rect 392176 329072 507860 329100
rect 392176 329060 392182 329072
rect 507854 329060 507860 329072
rect 507912 329060 507918 329112
rect 282914 328244 282920 328296
rect 282972 328284 282978 328296
rect 283190 328284 283196 328296
rect 282972 328256 283196 328284
rect 282972 328244 282978 328256
rect 283190 328244 283196 328256
rect 283248 328244 283254 328296
rect 318978 328176 318984 328228
rect 319036 328216 319042 328228
rect 319898 328216 319904 328228
rect 319036 328188 319904 328216
rect 319036 328176 319042 328188
rect 319898 328176 319904 328188
rect 319956 328176 319962 328228
rect 215294 327768 215300 327820
rect 215352 327808 215358 327820
rect 301314 327808 301320 327820
rect 215352 327780 301320 327808
rect 215352 327768 215358 327780
rect 301314 327768 301320 327780
rect 301372 327768 301378 327820
rect 346486 327768 346492 327820
rect 346544 327808 346550 327820
rect 347406 327808 347412 327820
rect 346544 327780 347412 327808
rect 346544 327768 346550 327780
rect 347406 327768 347412 327780
rect 347464 327768 347470 327820
rect 125594 327700 125600 327752
rect 125652 327740 125658 327752
rect 273438 327740 273444 327752
rect 125652 327712 273444 327740
rect 125652 327700 125658 327712
rect 273438 327700 273444 327712
rect 273496 327700 273502 327752
rect 394050 327700 394056 327752
rect 394108 327740 394114 327752
rect 514754 327740 514760 327752
rect 394108 327712 514760 327740
rect 394108 327700 394114 327712
rect 514754 327700 514760 327712
rect 514812 327700 514818 327752
rect 365714 327632 365720 327684
rect 365772 327672 365778 327684
rect 366358 327672 366364 327684
rect 365772 327644 366364 327672
rect 365772 327632 365778 327644
rect 366358 327632 366364 327644
rect 366416 327632 366422 327684
rect 393314 327564 393320 327616
rect 393372 327604 393378 327616
rect 393682 327604 393688 327616
rect 393372 327576 393688 327604
rect 393372 327564 393378 327576
rect 393682 327564 393688 327576
rect 393740 327564 393746 327616
rect 332686 327496 332692 327548
rect 332744 327536 332750 327548
rect 333054 327536 333060 327548
rect 332744 327508 333060 327536
rect 332744 327496 332750 327508
rect 333054 327496 333060 327508
rect 333112 327496 333118 327548
rect 283006 326884 283012 326936
rect 283064 326924 283070 326936
rect 283742 326924 283748 326936
rect 283064 326896 283748 326924
rect 283064 326884 283070 326896
rect 283742 326884 283748 326896
rect 283800 326884 283806 326936
rect 378318 326680 378324 326732
rect 378376 326680 378382 326732
rect 378336 326528 378364 326680
rect 280430 326476 280436 326528
rect 280488 326516 280494 326528
rect 280614 326516 280620 326528
rect 280488 326488 280620 326516
rect 280488 326476 280494 326488
rect 280614 326476 280620 326488
rect 280672 326476 280678 326528
rect 354950 326476 354956 326528
rect 355008 326516 355014 326528
rect 355134 326516 355140 326528
rect 355008 326488 355140 326516
rect 355008 326476 355014 326488
rect 355134 326476 355140 326488
rect 355192 326476 355198 326528
rect 375558 326476 375564 326528
rect 375616 326516 375622 326528
rect 375742 326516 375748 326528
rect 375616 326488 375748 326516
rect 375616 326476 375622 326488
rect 375742 326476 375748 326488
rect 375800 326476 375806 326528
rect 378318 326476 378324 326528
rect 378376 326476 378382 326528
rect 410058 326476 410064 326528
rect 410116 326516 410122 326528
rect 410334 326516 410340 326528
rect 410116 326488 410340 326516
rect 410116 326476 410122 326488
rect 410334 326476 410340 326488
rect 410392 326476 410398 326528
rect 193214 326408 193220 326460
rect 193272 326448 193278 326460
rect 293218 326448 293224 326460
rect 193272 326420 293224 326448
rect 193272 326408 193278 326420
rect 293218 326408 293224 326420
rect 293276 326408 293282 326460
rect 295518 326408 295524 326460
rect 295576 326408 295582 326460
rect 323026 326408 323032 326460
rect 323084 326448 323090 326460
rect 323946 326448 323952 326460
rect 323084 326420 323952 326448
rect 323084 326408 323090 326420
rect 323946 326408 323952 326420
rect 324004 326408 324010 326460
rect 328454 326408 328460 326460
rect 328512 326448 328518 326460
rect 329098 326448 329104 326460
rect 328512 326420 329104 326448
rect 328512 326408 328518 326420
rect 329098 326408 329104 326420
rect 329156 326408 329162 326460
rect 354674 326408 354680 326460
rect 354732 326448 354738 326460
rect 355686 326448 355692 326460
rect 354732 326420 355692 326448
rect 354732 326408 354738 326420
rect 355686 326408 355692 326420
rect 355744 326408 355750 326460
rect 356238 326408 356244 326460
rect 356296 326448 356302 326460
rect 356422 326448 356428 326460
rect 356296 326420 356428 326448
rect 356296 326408 356302 326420
rect 356422 326408 356428 326420
rect 356480 326408 356486 326460
rect 371234 326408 371240 326460
rect 371292 326448 371298 326460
rect 371786 326448 371792 326460
rect 371292 326420 371792 326448
rect 371292 326408 371298 326420
rect 371786 326408 371792 326420
rect 371844 326408 371850 326460
rect 372614 326408 372620 326460
rect 372672 326448 372678 326460
rect 373626 326448 373632 326460
rect 372672 326420 373632 326448
rect 372672 326408 372678 326420
rect 373626 326408 373632 326420
rect 373684 326408 373690 326460
rect 374178 326408 374184 326460
rect 374236 326448 374242 326460
rect 374730 326448 374736 326460
rect 374236 326420 374736 326448
rect 374236 326408 374242 326420
rect 374730 326408 374736 326420
rect 374788 326408 374794 326460
rect 375374 326408 375380 326460
rect 375432 326448 375438 326460
rect 376202 326448 376208 326460
rect 375432 326420 376208 326448
rect 375432 326408 375438 326420
rect 376202 326408 376208 326420
rect 376260 326408 376266 326460
rect 376846 326408 376852 326460
rect 376904 326448 376910 326460
rect 377674 326448 377680 326460
rect 376904 326420 377680 326448
rect 376904 326408 376910 326420
rect 377674 326408 377680 326420
rect 377732 326408 377738 326460
rect 378226 326408 378232 326460
rect 378284 326448 378290 326460
rect 379146 326448 379152 326460
rect 378284 326420 379152 326448
rect 378284 326408 378290 326420
rect 379146 326408 379152 326420
rect 379204 326408 379210 326460
rect 379514 326408 379520 326460
rect 379572 326448 379578 326460
rect 380526 326448 380532 326460
rect 379572 326420 380532 326448
rect 379572 326408 379578 326420
rect 380526 326408 380532 326420
rect 380584 326408 380590 326460
rect 381078 326408 381084 326460
rect 381136 326448 381142 326460
rect 381262 326448 381268 326460
rect 381136 326420 381268 326448
rect 381136 326408 381142 326420
rect 381262 326408 381268 326420
rect 381320 326408 381326 326460
rect 382274 326408 382280 326460
rect 382332 326448 382338 326460
rect 382734 326448 382740 326460
rect 382332 326420 382740 326448
rect 382332 326408 382338 326420
rect 382734 326408 382740 326420
rect 382792 326408 382798 326460
rect 383746 326408 383752 326460
rect 383804 326448 383810 326460
rect 384574 326448 384580 326460
rect 383804 326420 384580 326448
rect 383804 326408 383810 326420
rect 384574 326408 384580 326420
rect 384632 326408 384638 326460
rect 385218 326408 385224 326460
rect 385276 326448 385282 326460
rect 385678 326448 385684 326460
rect 385276 326420 385684 326448
rect 385276 326408 385282 326420
rect 385678 326408 385684 326420
rect 385736 326408 385742 326460
rect 386506 326408 386512 326460
rect 386564 326448 386570 326460
rect 387150 326448 387156 326460
rect 386564 326420 387156 326448
rect 386564 326408 386570 326420
rect 387150 326408 387156 326420
rect 387208 326408 387214 326460
rect 387794 326408 387800 326460
rect 387852 326448 387858 326460
rect 388622 326448 388628 326460
rect 387852 326420 388628 326448
rect 387852 326408 387858 326420
rect 388622 326408 388628 326420
rect 388680 326408 388686 326460
rect 398926 326408 398932 326460
rect 398984 326448 398990 326460
rect 399110 326448 399116 326460
rect 398984 326420 399116 326448
rect 398984 326408 398990 326420
rect 399110 326408 399116 326420
rect 399168 326408 399174 326460
rect 401686 326408 401692 326460
rect 401744 326448 401750 326460
rect 402514 326448 402520 326460
rect 401744 326420 402520 326448
rect 401744 326408 401750 326420
rect 402514 326408 402520 326420
rect 402572 326408 402578 326460
rect 403066 326408 403072 326460
rect 403124 326448 403130 326460
rect 403894 326448 403900 326460
rect 403124 326420 403900 326448
rect 403124 326408 403130 326420
rect 403894 326408 403900 326420
rect 403952 326408 403958 326460
rect 404446 326408 404452 326460
rect 404504 326448 404510 326460
rect 404630 326448 404636 326460
rect 404504 326420 404636 326448
rect 404504 326408 404510 326420
rect 404630 326408 404636 326420
rect 404688 326408 404694 326460
rect 405918 326408 405924 326460
rect 405976 326448 405982 326460
rect 406470 326448 406476 326460
rect 405976 326420 406476 326448
rect 405976 326408 405982 326420
rect 406470 326408 406476 326420
rect 406528 326408 406534 326460
rect 407114 326408 407120 326460
rect 407172 326448 407178 326460
rect 407574 326448 407580 326460
rect 407172 326420 407580 326448
rect 407172 326408 407178 326420
rect 407574 326408 407580 326420
rect 407632 326408 407638 326460
rect 409874 326408 409880 326460
rect 409932 326448 409938 326460
rect 410518 326448 410524 326460
rect 409932 326420 410524 326448
rect 409932 326408 409938 326420
rect 410518 326408 410524 326420
rect 410576 326408 410582 326460
rect 411346 326408 411352 326460
rect 411404 326448 411410 326460
rect 412358 326448 412364 326460
rect 411404 326420 412364 326448
rect 411404 326408 411410 326420
rect 412358 326408 412364 326420
rect 412416 326408 412422 326460
rect 4798 326340 4804 326392
rect 4856 326380 4862 326392
rect 234798 326380 234804 326392
rect 4856 326352 234804 326380
rect 4856 326340 4862 326352
rect 234798 326340 234804 326352
rect 234856 326340 234862 326392
rect 244274 326340 244280 326392
rect 244332 326380 244338 326392
rect 244734 326380 244740 326392
rect 244332 326352 244740 326380
rect 244332 326340 244338 326352
rect 244734 326340 244740 326352
rect 244792 326340 244798 326392
rect 245746 326340 245752 326392
rect 245804 326380 245810 326392
rect 246574 326380 246580 326392
rect 245804 326352 246580 326380
rect 245804 326340 245810 326352
rect 246574 326340 246580 326352
rect 246632 326340 246638 326392
rect 247034 326340 247040 326392
rect 247092 326380 247098 326392
rect 247954 326380 247960 326392
rect 247092 326352 247960 326380
rect 247092 326340 247098 326352
rect 247954 326340 247960 326352
rect 248012 326340 248018 326392
rect 249794 326340 249800 326392
rect 249852 326380 249858 326392
rect 250162 326380 250168 326392
rect 249852 326352 250168 326380
rect 249852 326340 249858 326352
rect 250162 326340 250168 326352
rect 250220 326340 250226 326392
rect 251174 326340 251180 326392
rect 251232 326380 251238 326392
rect 252002 326380 252008 326392
rect 251232 326352 252008 326380
rect 251232 326340 251238 326352
rect 252002 326340 252008 326352
rect 252060 326340 252066 326392
rect 273346 326340 273352 326392
rect 273404 326380 273410 326392
rect 274266 326380 274272 326392
rect 273404 326352 274272 326380
rect 273404 326340 273410 326352
rect 274266 326340 274272 326352
rect 274324 326340 274330 326392
rect 274634 326340 274640 326392
rect 274692 326380 274698 326392
rect 275002 326380 275008 326392
rect 274692 326352 275008 326380
rect 274692 326340 274698 326352
rect 275002 326340 275008 326352
rect 275060 326340 275066 326392
rect 276014 326340 276020 326392
rect 276072 326380 276078 326392
rect 276474 326380 276480 326392
rect 276072 326352 276480 326380
rect 276072 326340 276078 326352
rect 276474 326340 276480 326352
rect 276532 326340 276538 326392
rect 277486 326340 277492 326392
rect 277544 326380 277550 326392
rect 278314 326380 278320 326392
rect 277544 326352 278320 326380
rect 277544 326340 277550 326352
rect 278314 326340 278320 326352
rect 278372 326340 278378 326392
rect 278958 326340 278964 326392
rect 279016 326380 279022 326392
rect 279418 326380 279424 326392
rect 279016 326352 279424 326380
rect 279016 326340 279022 326352
rect 279418 326340 279424 326352
rect 279476 326340 279482 326392
rect 280246 326340 280252 326392
rect 280304 326380 280310 326392
rect 281258 326380 281264 326392
rect 280304 326352 281264 326380
rect 280304 326340 280310 326352
rect 281258 326340 281264 326352
rect 281316 326340 281322 326392
rect 281534 326340 281540 326392
rect 281592 326380 281598 326392
rect 281994 326380 282000 326392
rect 281592 326352 282000 326380
rect 281592 326340 281598 326352
rect 281994 326340 282000 326352
rect 282052 326340 282058 326392
rect 294230 326340 294236 326392
rect 294288 326380 294294 326392
rect 295150 326380 295156 326392
rect 294288 326352 295156 326380
rect 294288 326340 294294 326352
rect 295150 326340 295156 326352
rect 295208 326340 295214 326392
rect 249886 326272 249892 326324
rect 249944 326312 249950 326324
rect 250898 326312 250904 326324
rect 249944 326284 250904 326312
rect 249944 326272 249950 326284
rect 250898 326272 250904 326284
rect 250956 326272 250962 326324
rect 278774 326272 278780 326324
rect 278832 326312 278838 326324
rect 279786 326312 279792 326324
rect 278832 326284 279792 326312
rect 278832 326272 278838 326284
rect 279786 326272 279792 326284
rect 279844 326272 279850 326324
rect 295536 326256 295564 326408
rect 296990 326340 296996 326392
rect 297048 326380 297054 326392
rect 297634 326380 297640 326392
rect 297048 326352 297640 326380
rect 297048 326340 297054 326352
rect 297634 326340 297640 326352
rect 297692 326340 297698 326392
rect 299566 326340 299572 326392
rect 299624 326380 299630 326392
rect 300578 326380 300584 326392
rect 299624 326352 300584 326380
rect 299624 326340 299630 326352
rect 300578 326340 300584 326352
rect 300636 326340 300642 326392
rect 300854 326340 300860 326392
rect 300912 326380 300918 326392
rect 301682 326380 301688 326392
rect 300912 326352 301688 326380
rect 300912 326340 300918 326352
rect 301682 326340 301688 326352
rect 301740 326340 301746 326392
rect 321646 326340 321652 326392
rect 321704 326380 321710 326392
rect 322474 326380 322480 326392
rect 321704 326352 322480 326380
rect 321704 326340 321710 326352
rect 322474 326340 322480 326352
rect 322532 326340 322538 326392
rect 322934 326340 322940 326392
rect 322992 326380 322998 326392
rect 323578 326380 323584 326392
rect 322992 326352 323584 326380
rect 322992 326340 322998 326352
rect 323578 326340 323584 326352
rect 323636 326340 323642 326392
rect 327258 326340 327264 326392
rect 327316 326380 327322 326392
rect 327994 326380 328000 326392
rect 327316 326352 328000 326380
rect 327316 326340 327322 326352
rect 327994 326340 328000 326352
rect 328052 326340 328058 326392
rect 328638 326340 328644 326392
rect 328696 326380 328702 326392
rect 329466 326380 329472 326392
rect 328696 326352 329472 326380
rect 328696 326340 328702 326352
rect 329466 326340 329472 326352
rect 329524 326340 329530 326392
rect 329926 326340 329932 326392
rect 329984 326380 329990 326392
rect 330570 326380 330576 326392
rect 329984 326352 330576 326380
rect 329984 326340 329990 326352
rect 330570 326340 330576 326352
rect 330628 326340 330634 326392
rect 350534 326340 350540 326392
rect 350592 326380 350598 326392
rect 351362 326380 351368 326392
rect 350592 326352 351368 326380
rect 350592 326340 350598 326352
rect 351362 326340 351368 326352
rect 351420 326340 351426 326392
rect 354766 326340 354772 326392
rect 354824 326380 354830 326392
rect 355318 326380 355324 326392
rect 354824 326352 355324 326380
rect 354824 326340 354830 326352
rect 355318 326340 355324 326352
rect 355376 326340 355382 326392
rect 356054 326340 356060 326392
rect 356112 326380 356118 326392
rect 357158 326380 357164 326392
rect 356112 326352 357164 326380
rect 356112 326340 356118 326352
rect 357158 326340 357164 326352
rect 357216 326340 357222 326392
rect 364610 326340 364616 326392
rect 364668 326380 364674 326392
rect 419534 326380 419540 326392
rect 364668 326352 419540 326380
rect 364668 326340 364674 326352
rect 419534 326340 419540 326352
rect 419592 326340 419598 326392
rect 385034 326272 385040 326324
rect 385092 326312 385098 326324
rect 386046 326312 386052 326324
rect 385092 326284 386052 326312
rect 385092 326272 385098 326284
rect 386046 326272 386052 326284
rect 386104 326272 386110 326324
rect 386598 326272 386604 326324
rect 386656 326312 386662 326324
rect 387518 326312 387524 326324
rect 386656 326284 387524 326312
rect 386656 326272 386662 326284
rect 387518 326272 387524 326284
rect 387576 326272 387582 326324
rect 405734 326272 405740 326324
rect 405792 326312 405798 326324
rect 406838 326312 406844 326324
rect 405792 326284 406844 326312
rect 405792 326272 405798 326284
rect 406838 326272 406844 326284
rect 406896 326272 406902 326324
rect 295518 326204 295524 326256
rect 295576 326204 295582 326256
rect 410058 326204 410064 326256
rect 410116 326244 410122 326256
rect 410886 326244 410892 326256
rect 410116 326216 410892 326244
rect 410116 326204 410122 326216
rect 410886 326204 410892 326216
rect 410944 326204 410950 326256
rect 305270 326000 305276 326052
rect 305328 326040 305334 326052
rect 306098 326040 306104 326052
rect 305328 326012 306104 326040
rect 305328 326000 305334 326012
rect 306098 326000 306104 326012
rect 306156 326000 306162 326052
rect 371418 325728 371424 325780
rect 371476 325768 371482 325780
rect 372154 325768 372160 325780
rect 371476 325740 372160 325768
rect 371476 325728 371482 325740
rect 372154 325728 372160 325740
rect 372212 325728 372218 325780
rect 205634 325048 205640 325100
rect 205692 325088 205698 325100
rect 298278 325088 298284 325100
rect 205692 325060 298284 325088
rect 205692 325048 205698 325060
rect 298278 325048 298284 325060
rect 298336 325048 298342 325100
rect 164234 324980 164240 325032
rect 164292 325020 164298 325032
rect 276658 325020 276664 325032
rect 164292 324992 276664 325020
rect 164292 324980 164298 324992
rect 276658 324980 276664 324992
rect 276716 324980 276722 325032
rect 40034 324912 40040 324964
rect 40092 324952 40098 324964
rect 247310 324952 247316 324964
rect 40092 324924 247316 324952
rect 40092 324912 40098 324924
rect 247310 324912 247316 324924
rect 247368 324912 247374 324964
rect 363782 324912 363788 324964
rect 363840 324952 363846 324964
rect 416774 324952 416780 324964
rect 363840 324924 416780 324952
rect 363840 324912 363846 324924
rect 416774 324912 416780 324924
rect 416832 324912 416838 324964
rect 408494 324504 408500 324556
rect 408552 324544 408558 324556
rect 409046 324544 409052 324556
rect 408552 324516 409052 324544
rect 408552 324504 408558 324516
rect 409046 324504 409052 324516
rect 409104 324504 409110 324556
rect 407206 324232 407212 324284
rect 407264 324272 407270 324284
rect 407942 324272 407948 324284
rect 407264 324244 407948 324272
rect 407264 324232 407270 324244
rect 407942 324232 407948 324244
rect 408000 324232 408006 324284
rect 408586 323824 408592 323876
rect 408644 323864 408650 323876
rect 409414 323864 409420 323876
rect 408644 323836 409420 323864
rect 408644 323824 408650 323836
rect 409414 323824 409420 323836
rect 409472 323824 409478 323876
rect 128354 323620 128360 323672
rect 128412 323660 128418 323672
rect 274818 323660 274824 323672
rect 128412 323632 274824 323660
rect 128412 323620 128418 323632
rect 274818 323620 274824 323632
rect 274876 323620 274882 323672
rect 89714 323552 89720 323604
rect 89772 323592 89778 323604
rect 262582 323592 262588 323604
rect 89772 323564 262588 323592
rect 89772 323552 89778 323564
rect 262582 323552 262588 323564
rect 262640 323552 262646 323604
rect 280154 323552 280160 323604
rect 280212 323592 280218 323604
rect 280890 323592 280896 323604
rect 280212 323564 280896 323592
rect 280212 323552 280218 323564
rect 280890 323552 280896 323564
rect 280948 323552 280954 323604
rect 295426 323552 295432 323604
rect 295484 323592 295490 323604
rect 295610 323592 295616 323604
rect 295484 323564 295616 323592
rect 295484 323552 295490 323564
rect 295610 323552 295616 323564
rect 295668 323552 295674 323604
rect 325786 323552 325792 323604
rect 325844 323592 325850 323604
rect 325970 323592 325976 323604
rect 325844 323564 325976 323592
rect 325844 323552 325850 323564
rect 325970 323552 325976 323564
rect 326028 323552 326034 323604
rect 397730 323552 397736 323604
rect 397788 323592 397794 323604
rect 525794 323592 525800 323604
rect 397788 323564 525800 323592
rect 397788 323552 397794 323564
rect 525794 323552 525800 323564
rect 525852 323552 525858 323604
rect 358906 323212 358912 323264
rect 358964 323252 358970 323264
rect 359734 323252 359740 323264
rect 358964 323224 359740 323252
rect 358964 323212 358970 323224
rect 359734 323212 359740 323224
rect 359792 323212 359798 323264
rect 369854 323144 369860 323196
rect 369912 323184 369918 323196
rect 370682 323184 370688 323196
rect 369912 323156 370688 323184
rect 369912 323144 369918 323156
rect 370682 323144 370688 323156
rect 370740 323144 370746 323196
rect 380894 322736 380900 322788
rect 380952 322776 380958 322788
rect 381998 322776 382004 322788
rect 380952 322748 382004 322776
rect 380952 322736 380958 322748
rect 381998 322736 382004 322748
rect 382056 322736 382062 322788
rect 357618 322600 357624 322652
rect 357676 322640 357682 322652
rect 358262 322640 358268 322652
rect 357676 322612 358268 322640
rect 357676 322600 357682 322612
rect 358262 322600 358268 322612
rect 358320 322600 358326 322652
rect 358814 322532 358820 322584
rect 358872 322572 358878 322584
rect 359090 322572 359096 322584
rect 358872 322544 359096 322572
rect 358872 322532 358878 322544
rect 359090 322532 359096 322544
rect 359148 322532 359154 322584
rect 189074 322260 189080 322312
rect 189132 322300 189138 322312
rect 291930 322300 291936 322312
rect 189132 322272 291936 322300
rect 189132 322260 189138 322272
rect 291930 322260 291936 322272
rect 291988 322260 291994 322312
rect 51074 322192 51080 322244
rect 51132 322232 51138 322244
rect 250530 322232 250536 322244
rect 51132 322204 250536 322232
rect 51132 322192 51138 322204
rect 250530 322192 250536 322204
rect 250588 322192 250594 322244
rect 397638 322192 397644 322244
rect 397696 322232 397702 322244
rect 529934 322232 529940 322244
rect 397696 322204 529940 322232
rect 397696 322192 397702 322204
rect 529934 322192 529940 322204
rect 529992 322192 529998 322244
rect 387886 322124 387892 322176
rect 387944 322164 387950 322176
rect 388254 322164 388260 322176
rect 387944 322136 388260 322164
rect 387944 322124 387950 322136
rect 388254 322124 388260 322136
rect 388312 322124 388318 322176
rect 295334 322056 295340 322108
rect 295392 322096 295398 322108
rect 296162 322096 296168 322108
rect 295392 322068 296168 322096
rect 295392 322056 295398 322068
rect 296162 322056 296168 322068
rect 296220 322056 296226 322108
rect 329834 321580 329840 321632
rect 329892 321620 329898 321632
rect 330202 321620 330208 321632
rect 329892 321592 330208 321620
rect 329892 321580 329898 321592
rect 330202 321580 330208 321592
rect 330260 321580 330266 321632
rect 364886 320968 364892 321020
rect 364944 321008 364950 321020
rect 420914 321008 420920 321020
rect 364944 320980 420920 321008
rect 364944 320968 364950 320980
rect 420914 320968 420920 320980
rect 420972 320968 420978 321020
rect 385310 320900 385316 320952
rect 385368 320940 385374 320952
rect 487154 320940 487160 320952
rect 385368 320912 487160 320940
rect 385368 320900 385374 320912
rect 487154 320900 487160 320912
rect 487212 320900 487218 320952
rect 176654 320832 176660 320884
rect 176712 320872 176718 320884
rect 289906 320872 289912 320884
rect 176712 320844 289912 320872
rect 176712 320832 176718 320844
rect 289906 320832 289912 320844
rect 289964 320832 289970 320884
rect 292574 320832 292580 320884
rect 292632 320872 292638 320884
rect 292758 320872 292764 320884
rect 292632 320844 292764 320872
rect 292632 320832 292638 320844
rect 292758 320832 292764 320844
rect 292816 320832 292822 320884
rect 306374 320832 306380 320884
rect 306432 320872 306438 320884
rect 306558 320872 306564 320884
rect 306432 320844 306564 320872
rect 306432 320832 306438 320844
rect 306558 320832 306564 320844
rect 306616 320832 306622 320884
rect 413186 320832 413192 320884
rect 413244 320872 413250 320884
rect 576118 320872 576124 320884
rect 413244 320844 576124 320872
rect 413244 320832 413250 320844
rect 576118 320832 576124 320844
rect 576176 320832 576182 320884
rect 248414 320764 248420 320816
rect 248472 320804 248478 320816
rect 248598 320804 248604 320816
rect 248472 320776 248604 320804
rect 248472 320764 248478 320776
rect 248598 320764 248604 320776
rect 248656 320764 248662 320816
rect 3418 320084 3424 320136
rect 3476 320124 3482 320136
rect 232498 320124 232504 320136
rect 3476 320096 232504 320124
rect 3476 320084 3482 320096
rect 232498 320084 232504 320096
rect 232556 320084 232562 320136
rect 367370 319472 367376 319524
rect 367428 319512 367434 319524
rect 427814 319512 427820 319524
rect 367428 319484 427820 319512
rect 367428 319472 367434 319484
rect 427814 319472 427820 319484
rect 427872 319472 427878 319524
rect 223574 319404 223580 319456
rect 223632 319444 223638 319456
rect 303798 319444 303804 319456
rect 223632 319416 303804 319444
rect 223632 319404 223638 319416
rect 303798 319404 303804 319416
rect 303856 319404 303862 319456
rect 386690 319404 386696 319456
rect 386748 319444 386754 319456
rect 489914 319444 489920 319456
rect 386748 319416 489920 319444
rect 386748 319404 386754 319416
rect 489914 319404 489920 319416
rect 489972 319404 489978 319456
rect 370314 318112 370320 318164
rect 370372 318152 370378 318164
rect 438854 318152 438860 318164
rect 370372 318124 438860 318152
rect 370372 318112 370378 318124
rect 438854 318112 438860 318124
rect 438912 318112 438918 318164
rect 226334 318044 226340 318096
rect 226392 318084 226398 318096
rect 305178 318084 305184 318096
rect 226392 318056 305184 318084
rect 226392 318044 226398 318056
rect 305178 318044 305184 318056
rect 305236 318044 305242 318096
rect 386598 318044 386604 318096
rect 386656 318084 386662 318096
rect 494054 318084 494060 318096
rect 386656 318056 494060 318084
rect 386656 318044 386662 318056
rect 494054 318044 494060 318056
rect 494112 318044 494118 318096
rect 122834 316684 122840 316736
rect 122892 316724 122898 316736
rect 271966 316724 271972 316736
rect 122892 316696 271972 316724
rect 122892 316684 122898 316696
rect 271966 316684 271972 316696
rect 272024 316684 272030 316736
rect 387794 316684 387800 316736
rect 387852 316724 387858 316736
rect 498194 316724 498200 316736
rect 387852 316696 498200 316724
rect 387852 316684 387858 316696
rect 498194 316684 498200 316696
rect 498252 316684 498258 316736
rect 394694 315256 394700 315308
rect 394752 315296 394758 315308
rect 518894 315296 518900 315308
rect 394752 315268 518900 315296
rect 394752 315256 394758 315268
rect 518894 315256 518900 315268
rect 518952 315256 518958 315308
rect 391934 313896 391940 313948
rect 391992 313936 391998 313948
rect 511994 313936 512000 313948
rect 391992 313908 512000 313936
rect 391992 313896 391998 313908
rect 511994 313896 512000 313908
rect 512052 313896 512058 313948
rect 171134 312604 171140 312656
rect 171192 312644 171198 312656
rect 286410 312644 286416 312656
rect 171192 312616 286416 312644
rect 171192 312604 171198 312616
rect 286410 312604 286416 312616
rect 286468 312604 286474 312656
rect 64874 312536 64880 312588
rect 64932 312576 64938 312588
rect 254118 312576 254124 312588
rect 64932 312548 254124 312576
rect 64932 312536 64938 312548
rect 254118 312536 254124 312548
rect 254176 312536 254182 312588
rect 368750 312536 368756 312588
rect 368808 312576 368814 312588
rect 434714 312576 434720 312588
rect 368808 312548 434720 312576
rect 368808 312536 368814 312548
rect 434714 312536 434720 312548
rect 434772 312536 434778 312588
rect 400858 311108 400864 311160
rect 400916 311148 400922 311160
rect 532694 311148 532700 311160
rect 400916 311120 532700 311148
rect 400916 311108 400922 311120
rect 532694 311108 532700 311120
rect 532752 311108 532758 311160
rect 135254 309816 135260 309868
rect 135312 309856 135318 309868
rect 276198 309856 276204 309868
rect 135312 309828 276204 309856
rect 135312 309816 135318 309828
rect 276198 309816 276204 309828
rect 276256 309816 276262 309868
rect 81434 309748 81440 309800
rect 81492 309788 81498 309800
rect 259730 309788 259736 309800
rect 81492 309760 259736 309788
rect 81492 309748 81498 309760
rect 259730 309748 259736 309760
rect 259788 309748 259794 309800
rect 406010 309748 406016 309800
rect 406068 309788 406074 309800
rect 554774 309788 554780 309800
rect 406068 309760 554780 309788
rect 406068 309748 406074 309760
rect 554774 309748 554780 309760
rect 554832 309748 554838 309800
rect 132494 308456 132500 308508
rect 132552 308496 132558 308508
rect 274818 308496 274824 308508
rect 132552 308468 274824 308496
rect 132552 308456 132558 308468
rect 274818 308456 274824 308468
rect 274876 308456 274882 308508
rect 74534 308388 74540 308440
rect 74592 308428 74598 308440
rect 258350 308428 258356 308440
rect 74592 308400 258356 308428
rect 74592 308388 74598 308400
rect 258350 308388 258356 308400
rect 258408 308388 258414 308440
rect 408586 308388 408592 308440
rect 408644 308428 408650 308440
rect 564434 308428 564440 308440
rect 408644 308400 564440 308428
rect 408644 308388 408650 308400
rect 564434 308388 564440 308400
rect 564492 308388 564498 308440
rect 207014 307096 207020 307148
rect 207072 307136 207078 307148
rect 294598 307136 294604 307148
rect 207072 307108 294604 307136
rect 207072 307096 207078 307108
rect 294598 307096 294604 307108
rect 294656 307096 294662 307148
rect 60734 307028 60740 307080
rect 60792 307068 60798 307080
rect 253198 307068 253204 307080
rect 60792 307040 253204 307068
rect 60792 307028 60798 307040
rect 253198 307028 253204 307040
rect 253256 307028 253262 307080
rect 409874 307028 409880 307080
rect 409932 307068 409938 307080
rect 568574 307068 568580 307080
rect 409932 307040 568580 307068
rect 409932 307028 409938 307040
rect 568574 307028 568580 307040
rect 568632 307028 568638 307080
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 383010 306320 383016 306332
rect 3384 306292 383016 306320
rect 3384 306280 3390 306292
rect 383010 306280 383016 306292
rect 383068 306280 383074 306332
rect 371510 305668 371516 305720
rect 371568 305708 371574 305720
rect 441614 305708 441620 305720
rect 371568 305680 441620 305708
rect 371568 305668 371574 305680
rect 441614 305668 441620 305680
rect 441672 305668 441678 305720
rect 390830 305600 390836 305652
rect 390888 305640 390894 305652
rect 505094 305640 505100 305652
rect 390888 305612 505100 305640
rect 390888 305600 390894 305612
rect 505094 305600 505100 305612
rect 505152 305600 505158 305652
rect 209774 304308 209780 304360
rect 209832 304348 209838 304360
rect 297450 304348 297456 304360
rect 209832 304320 297456 304348
rect 209832 304308 209838 304320
rect 297450 304308 297456 304320
rect 297508 304308 297514 304360
rect 53834 304240 53840 304292
rect 53892 304280 53898 304292
rect 251358 304280 251364 304292
rect 53892 304252 251364 304280
rect 53892 304240 53898 304252
rect 251358 304240 251364 304252
rect 251416 304240 251422 304292
rect 379606 304240 379612 304292
rect 379664 304280 379670 304292
rect 470594 304280 470600 304292
rect 379664 304252 470600 304280
rect 379664 304240 379670 304252
rect 470594 304240 470600 304252
rect 470652 304240 470658 304292
rect 157334 302948 157340 303000
rect 157392 302988 157398 303000
rect 283190 302988 283196 303000
rect 157392 302960 283196 302988
rect 157392 302948 157398 302960
rect 283190 302948 283196 302960
rect 283248 302948 283254 303000
rect 25498 302880 25504 302932
rect 25556 302920 25562 302932
rect 241790 302920 241796 302932
rect 25556 302892 241796 302920
rect 25556 302880 25562 302892
rect 241790 302880 241796 302892
rect 241848 302880 241854 302932
rect 146294 301452 146300 301504
rect 146352 301492 146358 301504
rect 280430 301492 280436 301504
rect 146352 301464 280436 301492
rect 146352 301452 146358 301464
rect 280430 301452 280436 301464
rect 280488 301452 280494 301504
rect 393498 301452 393504 301504
rect 393556 301492 393562 301504
rect 513374 301492 513380 301504
rect 393556 301464 513380 301492
rect 393556 301452 393562 301464
rect 513374 301452 513380 301464
rect 513432 301452 513438 301504
rect 143534 300092 143540 300144
rect 143592 300132 143598 300144
rect 279050 300132 279056 300144
rect 143592 300104 279056 300132
rect 143592 300092 143598 300104
rect 279050 300092 279056 300104
rect 279108 300092 279114 300144
rect 397546 300092 397552 300144
rect 397604 300132 397610 300144
rect 527174 300132 527180 300144
rect 397604 300104 527180 300132
rect 397604 300092 397610 300104
rect 527174 300092 527180 300104
rect 527232 300092 527238 300144
rect 424318 299412 424324 299464
rect 424376 299452 424382 299464
rect 580166 299452 580172 299464
rect 424376 299424 580172 299452
rect 424376 299412 424382 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 365898 298732 365904 298784
rect 365956 298772 365962 298784
rect 423766 298772 423772 298784
rect 365956 298744 423772 298772
rect 365956 298732 365962 298744
rect 423766 298732 423772 298744
rect 423824 298732 423830 298784
rect 400306 297372 400312 297424
rect 400364 297412 400370 297424
rect 536834 297412 536840 297424
rect 400364 297384 536840 297412
rect 400364 297372 400370 297384
rect 536834 297372 536840 297384
rect 536892 297372 536898 297424
rect 403066 295944 403072 295996
rect 403124 295984 403130 295996
rect 547874 295984 547880 295996
rect 403124 295956 547880 295984
rect 403124 295944 403130 295956
rect 547874 295944 547880 295956
rect 547932 295944 547938 295996
rect 407298 294584 407304 294636
rect 407356 294624 407362 294636
rect 557534 294624 557540 294636
rect 407356 294596 557540 294624
rect 407356 294584 407362 294596
rect 557534 294584 557540 294596
rect 557592 294584 557598 294636
rect 2866 293904 2872 293956
rect 2924 293944 2930 293956
rect 10318 293944 10324 293956
rect 2924 293916 10324 293944
rect 2924 293904 2930 293916
rect 10318 293904 10324 293916
rect 10376 293904 10382 293956
rect 413278 293224 413284 293276
rect 413336 293264 413342 293276
rect 572806 293264 572812 293276
rect 413336 293236 572812 293264
rect 413336 293224 413342 293236
rect 572806 293224 572812 293236
rect 572864 293224 572870 293276
rect 147674 291796 147680 291848
rect 147732 291836 147738 291848
rect 280338 291836 280344 291848
rect 147732 291808 280344 291836
rect 147732 291796 147738 291808
rect 280338 291796 280344 291808
rect 280396 291796 280402 291848
rect 398926 291796 398932 291848
rect 398984 291836 398990 291848
rect 531314 291836 531320 291848
rect 398984 291808 531320 291836
rect 398984 291796 398990 291808
rect 531314 291796 531320 291808
rect 531372 291796 531378 291848
rect 136634 290436 136640 290488
rect 136692 290476 136698 290488
rect 277578 290476 277584 290488
rect 136692 290448 277584 290476
rect 136692 290436 136698 290448
rect 277578 290436 277584 290448
rect 277636 290436 277642 290488
rect 402974 290436 402980 290488
rect 403032 290476 403038 290488
rect 545114 290476 545120 290488
rect 403032 290448 545120 290476
rect 403032 290436 403038 290448
rect 545114 290436 545120 290448
rect 545172 290436 545178 290488
rect 179414 289144 179420 289196
rect 179472 289184 179478 289196
rect 287698 289184 287704 289196
rect 179472 289156 287704 289184
rect 179472 289144 179478 289156
rect 287698 289144 287704 289156
rect 287756 289144 287762 289196
rect 35894 289076 35900 289128
rect 35952 289116 35958 289128
rect 244918 289116 244924 289128
rect 35952 289088 244924 289116
rect 35952 289076 35958 289088
rect 244918 289076 244924 289088
rect 244976 289076 244982 289128
rect 405918 289076 405924 289128
rect 405976 289116 405982 289128
rect 556154 289116 556160 289128
rect 405976 289088 556160 289116
rect 405976 289076 405982 289088
rect 556154 289076 556160 289088
rect 556212 289076 556218 289128
rect 139394 287648 139400 287700
rect 139452 287688 139458 287700
rect 273898 287688 273904 287700
rect 139452 287660 273904 287688
rect 139452 287648 139458 287660
rect 273898 287648 273904 287660
rect 273956 287648 273962 287700
rect 411438 287648 411444 287700
rect 411496 287688 411502 287700
rect 571978 287688 571984 287700
rect 411496 287660 571984 287688
rect 411496 287648 411502 287660
rect 571978 287648 571984 287660
rect 572036 287648 572042 287700
rect 178034 286356 178040 286408
rect 178092 286396 178098 286408
rect 289170 286396 289176 286408
rect 178092 286368 289176 286396
rect 178092 286356 178098 286368
rect 289170 286356 289176 286368
rect 289228 286356 289234 286408
rect 354950 286356 354956 286408
rect 355008 286396 355014 286408
rect 387794 286396 387800 286408
rect 355008 286368 387800 286396
rect 355008 286356 355014 286368
rect 387794 286356 387800 286368
rect 387852 286356 387858 286408
rect 118694 286288 118700 286340
rect 118752 286328 118758 286340
rect 269758 286328 269764 286340
rect 118752 286300 269764 286328
rect 118752 286288 118758 286300
rect 269758 286288 269764 286300
rect 269816 286288 269822 286340
rect 378410 286288 378416 286340
rect 378468 286328 378474 286340
rect 465166 286328 465172 286340
rect 378468 286300 465172 286328
rect 378468 286288 378474 286300
rect 465166 286288 465172 286300
rect 465224 286288 465230 286340
rect 182174 284996 182180 285048
rect 182232 285036 182238 285048
rect 286318 285036 286324 285048
rect 182232 285008 286324 285036
rect 182232 284996 182238 285008
rect 286318 284996 286324 285008
rect 286376 284996 286382 285048
rect 356330 284996 356336 285048
rect 356388 285036 356394 285048
rect 394694 285036 394700 285048
rect 356388 285008 394700 285036
rect 356388 284996 356394 285008
rect 394694 284996 394700 285008
rect 394752 284996 394758 285048
rect 62114 284928 62120 284980
rect 62172 284968 62178 284980
rect 254026 284968 254032 284980
rect 62172 284940 254032 284968
rect 62172 284928 62178 284940
rect 254026 284928 254032 284940
rect 254084 284928 254090 284980
rect 285674 284928 285680 284980
rect 285732 284968 285738 284980
rect 323210 284968 323216 284980
rect 285732 284940 323216 284968
rect 285732 284928 285738 284940
rect 323210 284928 323216 284940
rect 323268 284928 323274 284980
rect 381078 284928 381084 284980
rect 381136 284968 381142 284980
rect 473354 284968 473360 284980
rect 381136 284940 473360 284968
rect 381136 284928 381142 284940
rect 473354 284928 473360 284940
rect 473412 284928 473418 284980
rect 184934 283636 184940 283688
rect 184992 283676 184998 283688
rect 291378 283676 291384 283688
rect 184992 283648 291384 283676
rect 184992 283636 184998 283648
rect 291378 283636 291384 283648
rect 291436 283636 291442 283688
rect 360470 283636 360476 283688
rect 360528 283676 360534 283688
rect 408586 283676 408592 283688
rect 360528 283648 408592 283676
rect 360528 283636 360534 283648
rect 408586 283636 408592 283648
rect 408644 283636 408650 283688
rect 10318 283568 10324 283620
rect 10376 283608 10382 283620
rect 236086 283608 236092 283620
rect 10376 283580 236092 283608
rect 10376 283568 10382 283580
rect 236086 283568 236092 283580
rect 236144 283568 236150 283620
rect 390738 283568 390744 283620
rect 390796 283608 390802 283620
rect 506474 283608 506480 283620
rect 390796 283580 506480 283608
rect 390796 283568 390802 283580
rect 506474 283568 506480 283580
rect 506532 283568 506538 283620
rect 195974 282208 195980 282260
rect 196032 282248 196038 282260
rect 295518 282248 295524 282260
rect 196032 282220 295524 282248
rect 196032 282208 196038 282220
rect 295518 282208 295524 282220
rect 295576 282208 295582 282260
rect 363138 282208 363144 282260
rect 363196 282248 363202 282260
rect 415394 282248 415400 282260
rect 363196 282220 415400 282248
rect 363196 282208 363202 282220
rect 415394 282208 415400 282220
rect 415452 282208 415458 282260
rect 121454 282140 121460 282192
rect 121512 282180 121518 282192
rect 271138 282180 271144 282192
rect 121512 282152 271144 282180
rect 121512 282140 121518 282152
rect 271138 282140 271144 282152
rect 271196 282140 271202 282192
rect 394878 282140 394884 282192
rect 394936 282180 394942 282192
rect 520274 282180 520280 282192
rect 394936 282152 520280 282180
rect 394936 282140 394942 282152
rect 520274 282140 520280 282152
rect 520332 282140 520338 282192
rect 200114 280848 200120 280900
rect 200172 280888 200178 280900
rect 295978 280888 295984 280900
rect 200172 280860 295984 280888
rect 200172 280848 200178 280860
rect 295978 280848 295984 280860
rect 296036 280848 296042 280900
rect 365806 280848 365812 280900
rect 365864 280888 365870 280900
rect 426434 280888 426440 280900
rect 365864 280860 426440 280888
rect 365864 280848 365870 280860
rect 426434 280848 426440 280860
rect 426492 280848 426498 280900
rect 16574 280780 16580 280832
rect 16632 280820 16638 280832
rect 239398 280820 239404 280832
rect 16632 280792 239404 280820
rect 16632 280780 16638 280792
rect 239398 280780 239404 280792
rect 239456 280780 239462 280832
rect 404538 280780 404544 280832
rect 404596 280820 404602 280832
rect 552014 280820 552020 280832
rect 404596 280792 552020 280820
rect 404596 280780 404602 280792
rect 552014 280780 552020 280792
rect 552072 280780 552078 280832
rect 296714 279624 296720 279676
rect 296772 279664 296778 279676
rect 322198 279664 322204 279676
rect 296772 279636 322204 279664
rect 296772 279624 296778 279636
rect 322198 279624 322204 279636
rect 322256 279624 322262 279676
rect 202874 279488 202880 279540
rect 202932 279528 202938 279540
rect 296990 279528 296996 279540
rect 202932 279500 296996 279528
rect 202932 279488 202938 279500
rect 296990 279488 296996 279500
rect 297048 279488 297054 279540
rect 103514 279420 103520 279472
rect 103572 279460 103578 279472
rect 264238 279460 264244 279472
rect 103572 279432 264244 279460
rect 103572 279420 103578 279432
rect 264238 279420 264244 279432
rect 264296 279420 264302 279472
rect 372798 279420 372804 279472
rect 372856 279460 372862 279472
rect 448514 279460 448520 279472
rect 372856 279432 448520 279460
rect 372856 279420 372862 279432
rect 448514 279420 448520 279432
rect 448572 279420 448578 279472
rect 213914 278060 213920 278112
rect 213972 278100 213978 278112
rect 300946 278100 300952 278112
rect 213972 278072 300952 278100
rect 213972 278060 213978 278072
rect 300946 278060 300952 278072
rect 301004 278060 301010 278112
rect 85574 277992 85580 278044
rect 85632 278032 85638 278044
rect 261110 278032 261116 278044
rect 85632 278004 261116 278032
rect 85632 277992 85638 278004
rect 261110 277992 261116 278004
rect 261168 277992 261174 278044
rect 374270 277992 374276 278044
rect 374328 278032 374334 278044
rect 451274 278032 451280 278044
rect 374328 278004 451280 278032
rect 374328 277992 374334 278004
rect 451274 277992 451280 278004
rect 451332 277992 451338 278044
rect 220814 276700 220820 276752
rect 220872 276740 220878 276752
rect 302326 276740 302332 276752
rect 220872 276712 302332 276740
rect 220872 276700 220878 276712
rect 302326 276700 302332 276712
rect 302384 276700 302390 276752
rect 69014 276632 69020 276684
rect 69072 276672 69078 276684
rect 255590 276672 255596 276684
rect 69072 276644 255596 276672
rect 69072 276632 69078 276644
rect 255590 276632 255596 276644
rect 255648 276632 255654 276684
rect 375558 276632 375564 276684
rect 375616 276672 375622 276684
rect 455414 276672 455420 276684
rect 375616 276644 455420 276672
rect 375616 276632 375622 276644
rect 455414 276632 455420 276644
rect 455472 276632 455478 276684
rect 231854 275340 231860 275392
rect 231912 275380 231918 275392
rect 306558 275380 306564 275392
rect 231912 275352 306564 275380
rect 231912 275340 231918 275352
rect 306558 275340 306564 275352
rect 306616 275340 306622 275392
rect 11698 275272 11704 275324
rect 11756 275312 11762 275324
rect 234706 275312 234712 275324
rect 11756 275284 234712 275312
rect 11756 275272 11762 275284
rect 234706 275272 234712 275284
rect 234764 275272 234770 275324
rect 376938 275272 376944 275324
rect 376996 275312 377002 275324
rect 458174 275312 458180 275324
rect 376996 275284 458180 275312
rect 376996 275272 377002 275284
rect 458174 275272 458180 275284
rect 458232 275272 458238 275324
rect 274818 274048 274824 274100
rect 274876 274088 274882 274100
rect 319070 274088 319076 274100
rect 274876 274060 319076 274088
rect 274876 274048 274882 274060
rect 319070 274048 319076 274060
rect 319128 274048 319134 274100
rect 129734 273912 129740 273964
rect 129792 273952 129798 273964
rect 274634 273952 274640 273964
rect 129792 273924 274640 273952
rect 129792 273912 129798 273924
rect 274634 273912 274640 273924
rect 274692 273912 274698 273964
rect 376846 273912 376852 273964
rect 376904 273952 376910 273964
rect 462314 273952 462320 273964
rect 376904 273924 462320 273952
rect 376904 273912 376910 273924
rect 462314 273912 462320 273924
rect 462372 273912 462378 273964
rect 460198 273164 460204 273216
rect 460256 273204 460262 273216
rect 580166 273204 580172 273216
rect 460256 273176 580172 273204
rect 460256 273164 460262 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 150434 272484 150440 272536
rect 150492 272524 150498 272536
rect 280246 272524 280252 272536
rect 150492 272496 280252 272524
rect 150492 272484 150498 272496
rect 280246 272484 280252 272496
rect 280304 272484 280310 272536
rect 359090 272484 359096 272536
rect 359148 272524 359154 272536
rect 402974 272524 402980 272536
rect 359148 272496 402980 272524
rect 359148 272484 359154 272496
rect 402974 272484 402980 272496
rect 403032 272484 403038 272536
rect 153194 271124 153200 271176
rect 153252 271164 153258 271176
rect 281718 271164 281724 271176
rect 153252 271136 281724 271164
rect 153252 271124 153258 271136
rect 281718 271124 281724 271136
rect 281776 271124 281782 271176
rect 381538 271124 381544 271176
rect 381596 271164 381602 271176
rect 469214 271164 469220 271176
rect 381596 271136 469220 271164
rect 381596 271124 381602 271136
rect 469214 271124 469220 271136
rect 469272 271124 469278 271176
rect 161474 269764 161480 269816
rect 161532 269804 161538 269816
rect 284478 269804 284484 269816
rect 161532 269776 284484 269804
rect 161532 269764 161538 269776
rect 284478 269764 284484 269776
rect 284536 269764 284542 269816
rect 383838 269764 383844 269816
rect 383896 269804 383902 269816
rect 481634 269804 481640 269816
rect 383896 269776 481640 269804
rect 383896 269764 383902 269776
rect 481634 269764 481640 269776
rect 481692 269764 481698 269816
rect 165614 268336 165620 268388
rect 165672 268376 165678 268388
rect 285858 268376 285864 268388
rect 165672 268348 285864 268376
rect 165672 268336 165678 268348
rect 285858 268336 285864 268348
rect 285916 268336 285922 268388
rect 383746 268336 383752 268388
rect 383804 268376 383810 268388
rect 484394 268376 484400 268388
rect 383804 268348 484400 268376
rect 383804 268336 383810 268348
rect 484394 268336 484400 268348
rect 484452 268336 484458 268388
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 231118 267696 231124 267708
rect 3292 267668 231124 267696
rect 3292 267656 3298 267668
rect 231118 267656 231124 267668
rect 231176 267656 231182 267708
rect 222194 266976 222200 267028
rect 222252 267016 222258 267028
rect 303706 267016 303712 267028
rect 222252 266988 303712 267016
rect 222252 266976 222258 266988
rect 303706 266976 303712 266988
rect 303764 266976 303770 267028
rect 385218 266976 385224 267028
rect 385276 267016 385282 267028
rect 488534 267016 488540 267028
rect 385276 266988 488540 267016
rect 385276 266976 385282 266988
rect 488534 266976 488540 266988
rect 488592 266976 488598 267028
rect 168466 265616 168472 265668
rect 168524 265656 168530 265668
rect 287238 265656 287244 265668
rect 168524 265628 287244 265656
rect 168524 265616 168530 265628
rect 287238 265616 287244 265628
rect 287296 265616 287302 265668
rect 386414 265616 386420 265668
rect 386472 265656 386478 265668
rect 491294 265656 491300 265668
rect 386472 265628 491300 265656
rect 386472 265616 386478 265628
rect 491294 265616 491300 265628
rect 491352 265616 491358 265668
rect 172514 264188 172520 264240
rect 172572 264228 172578 264240
rect 287146 264228 287152 264240
rect 172572 264200 287152 264228
rect 172572 264188 172578 264200
rect 287146 264188 287152 264200
rect 287204 264188 287210 264240
rect 387978 264188 387984 264240
rect 388036 264228 388042 264240
rect 495434 264228 495440 264240
rect 388036 264200 495440 264228
rect 388036 264188 388042 264200
rect 495434 264188 495440 264200
rect 495492 264188 495498 264240
rect 183554 262828 183560 262880
rect 183612 262868 183618 262880
rect 291286 262868 291292 262880
rect 183612 262840 291292 262868
rect 183612 262828 183618 262840
rect 291286 262828 291292 262840
rect 291344 262828 291350 262880
rect 389174 262828 389180 262880
rect 389232 262868 389238 262880
rect 498286 262868 498292 262880
rect 389232 262840 498292 262868
rect 389232 262828 389238 262840
rect 498286 262828 498292 262840
rect 498344 262828 498350 262880
rect 292574 261536 292580 261588
rect 292632 261576 292638 261588
rect 324590 261576 324596 261588
rect 292632 261548 324596 261576
rect 292632 261536 292638 261548
rect 324590 261536 324596 261548
rect 324648 261536 324654 261588
rect 186314 261468 186320 261520
rect 186372 261508 186378 261520
rect 292758 261508 292764 261520
rect 186372 261480 292764 261508
rect 186372 261468 186378 261480
rect 292758 261468 292764 261480
rect 292816 261468 292822 261520
rect 354858 261468 354864 261520
rect 354916 261508 354922 261520
rect 389174 261508 389180 261520
rect 354916 261480 389180 261508
rect 354916 261468 354922 261480
rect 389174 261468 389180 261480
rect 389232 261468 389238 261520
rect 389358 261468 389364 261520
rect 389416 261508 389422 261520
rect 502334 261508 502340 261520
rect 389416 261480 502340 261508
rect 389416 261468 389422 261480
rect 502334 261468 502340 261480
rect 502392 261468 502398 261520
rect 190454 260108 190460 260160
rect 190512 260148 190518 260160
rect 292850 260148 292856 260160
rect 190512 260120 292856 260148
rect 190512 260108 190518 260120
rect 292850 260108 292856 260120
rect 292908 260108 292914 260160
rect 356238 260108 356244 260160
rect 356296 260148 356302 260160
rect 391934 260148 391940 260160
rect 356296 260120 391940 260148
rect 356296 260108 356302 260120
rect 391934 260108 391940 260120
rect 391992 260108 391998 260160
rect 392118 260108 392124 260160
rect 392176 260148 392182 260160
rect 509234 260148 509240 260160
rect 392176 260120 509240 260148
rect 392176 260108 392182 260120
rect 509234 260108 509240 260120
rect 509292 260108 509298 260160
rect 445018 259360 445024 259412
rect 445076 259400 445082 259412
rect 580166 259400 580172 259412
rect 445076 259372 580172 259400
rect 445076 259360 445082 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 193306 258680 193312 258732
rect 193364 258720 193370 258732
rect 294138 258720 294144 258732
rect 193364 258692 294144 258720
rect 193364 258680 193370 258692
rect 294138 258680 294144 258692
rect 294196 258680 294202 258732
rect 367278 258680 367284 258732
rect 367336 258720 367342 258732
rect 432046 258720 432052 258732
rect 367336 258692 432052 258720
rect 367336 258680 367342 258692
rect 432046 258680 432052 258692
rect 432104 258680 432110 258732
rect 197354 257320 197360 257372
rect 197412 257360 197418 257372
rect 295426 257360 295432 257372
rect 197412 257332 295432 257360
rect 197412 257320 197418 257332
rect 295426 257320 295432 257332
rect 295484 257320 295490 257372
rect 393406 257320 393412 257372
rect 393464 257360 393470 257372
rect 516134 257360 516140 257372
rect 393464 257332 516140 257360
rect 393464 257320 393470 257332
rect 516134 257320 516140 257332
rect 516192 257320 516198 257372
rect 204254 256028 204260 256080
rect 204312 256068 204318 256080
rect 298186 256068 298192 256080
rect 204312 256040 298192 256068
rect 204312 256028 204318 256040
rect 298186 256028 298192 256040
rect 298244 256028 298250 256080
rect 41414 255960 41420 256012
rect 41472 256000 41478 256012
rect 247218 256000 247224 256012
rect 41472 255972 247224 256000
rect 41472 255960 41478 255972
rect 247218 255960 247224 255972
rect 247276 255960 247282 256012
rect 357618 255960 357624 256012
rect 357676 256000 357682 256012
rect 398926 256000 398932 256012
rect 357676 255972 398932 256000
rect 357676 255960 357682 255972
rect 398926 255960 398932 255972
rect 398984 255960 398990 256012
rect 399018 255960 399024 256012
rect 399076 256000 399082 256012
rect 534074 256000 534080 256012
rect 399076 255972 534080 256000
rect 399076 255960 399082 255972
rect 534074 255960 534080 255972
rect 534132 255960 534138 256012
rect 3326 255212 3332 255264
rect 3384 255252 3390 255264
rect 17218 255252 17224 255264
rect 3384 255224 17224 255252
rect 3384 255212 3390 255224
rect 17218 255212 17224 255224
rect 17276 255212 17282 255264
rect 208394 254600 208400 254652
rect 208452 254640 208458 254652
rect 298370 254640 298376 254652
rect 208452 254612 298376 254640
rect 208452 254600 208458 254612
rect 298370 254600 298376 254612
rect 298428 254600 298434 254652
rect 34514 254532 34520 254584
rect 34572 254572 34578 254584
rect 245838 254572 245844 254584
rect 34572 254544 245844 254572
rect 34572 254532 34578 254544
rect 245838 254532 245844 254544
rect 245896 254532 245902 254584
rect 358998 254532 359004 254584
rect 359056 254572 359062 254584
rect 400306 254572 400312 254584
rect 359056 254544 400312 254572
rect 359056 254532 359062 254544
rect 400306 254532 400312 254544
rect 400364 254532 400370 254584
rect 400398 254532 400404 254584
rect 400456 254572 400462 254584
rect 538214 254572 538220 254584
rect 400456 254544 538220 254572
rect 400456 254532 400462 254544
rect 538214 254532 538220 254544
rect 538272 254532 538278 254584
rect 299474 253376 299480 253428
rect 299532 253416 299538 253428
rect 320818 253416 320824 253428
rect 299532 253388 320824 253416
rect 299532 253376 299538 253388
rect 320818 253376 320824 253388
rect 320876 253376 320882 253428
rect 211154 253240 211160 253292
rect 211212 253280 211218 253292
rect 299750 253280 299756 253292
rect 211212 253252 299756 253280
rect 211212 253240 211218 253252
rect 299750 253240 299756 253252
rect 299808 253240 299814 253292
rect 24118 253172 24124 253224
rect 24176 253212 24182 253224
rect 240318 253212 240324 253224
rect 24176 253184 240324 253212
rect 24176 253172 24182 253184
rect 240318 253172 240324 253184
rect 240376 253172 240382 253224
rect 404446 253172 404452 253224
rect 404504 253212 404510 253224
rect 547966 253212 547972 253224
rect 404504 253184 547972 253212
rect 404504 253172 404510 253184
rect 547966 253172 547972 253184
rect 548024 253172 548030 253224
rect 303614 252016 303620 252068
rect 303672 252056 303678 252068
rect 328730 252056 328736 252068
rect 303672 252028 328736 252056
rect 303672 252016 303678 252028
rect 328730 252016 328736 252028
rect 328788 252016 328794 252068
rect 226426 251880 226432 251932
rect 226484 251920 226490 251932
rect 303890 251920 303896 251932
rect 226484 251892 303896 251920
rect 226484 251880 226490 251892
rect 303890 251880 303896 251892
rect 303948 251880 303954 251932
rect 28994 251812 29000 251864
rect 29052 251852 29058 251864
rect 243078 251852 243084 251864
rect 29052 251824 243084 251852
rect 29052 251812 29058 251824
rect 243078 251812 243084 251824
rect 243136 251812 243142 251864
rect 408678 251812 408684 251864
rect 408736 251852 408742 251864
rect 563054 251852 563060 251864
rect 408736 251824 563060 251852
rect 408736 251812 408742 251824
rect 563054 251812 563060 251824
rect 563112 251812 563118 251864
rect 229094 250520 229100 250572
rect 229152 250560 229158 250572
rect 305086 250560 305092 250572
rect 229152 250532 305092 250560
rect 229152 250520 229158 250532
rect 305086 250520 305092 250532
rect 305144 250520 305150 250572
rect 20714 250452 20720 250504
rect 20772 250492 20778 250504
rect 241698 250492 241704 250504
rect 20772 250464 241704 250492
rect 20772 250452 20778 250464
rect 241698 250452 241704 250464
rect 241756 250452 241762 250504
rect 364978 250452 364984 250504
rect 365036 250492 365042 250504
rect 409874 250492 409880 250504
rect 365036 250464 409880 250492
rect 365036 250452 365042 250464
rect 409874 250452 409880 250464
rect 409932 250452 409938 250504
rect 410150 250452 410156 250504
rect 410208 250492 410214 250504
rect 565814 250492 565820 250504
rect 410208 250464 565820 250492
rect 410208 250452 410214 250464
rect 565814 250452 565820 250464
rect 565872 250452 565878 250504
rect 276198 249160 276204 249212
rect 276256 249200 276262 249212
rect 318978 249200 318984 249212
rect 276256 249172 318984 249200
rect 276256 249160 276262 249172
rect 318978 249160 318984 249172
rect 319036 249160 319042 249212
rect 133874 249024 133880 249076
rect 133932 249064 133938 249076
rect 276106 249064 276112 249076
rect 133932 249036 276112 249064
rect 133932 249024 133938 249036
rect 276106 249024 276112 249036
rect 276164 249024 276170 249076
rect 410058 249024 410064 249076
rect 410116 249064 410122 249076
rect 569954 249064 569960 249076
rect 410116 249036 569960 249064
rect 410116 249024 410122 249036
rect 569954 249024 569960 249036
rect 570012 249024 570018 249076
rect 233234 247732 233240 247784
rect 233292 247772 233298 247784
rect 306466 247772 306472 247784
rect 233292 247744 306472 247772
rect 233292 247732 233298 247744
rect 306466 247732 306472 247744
rect 306524 247732 306530 247784
rect 6914 247664 6920 247716
rect 6972 247704 6978 247716
rect 233970 247704 233976 247716
rect 6972 247676 233976 247704
rect 6972 247664 6978 247676
rect 233970 247664 233976 247676
rect 234028 247664 234034 247716
rect 385126 247664 385132 247716
rect 385184 247704 385190 247716
rect 485774 247704 485780 247716
rect 385184 247676 485780 247704
rect 385184 247664 385190 247676
rect 485774 247664 485780 247676
rect 485832 247664 485838 247716
rect 386506 246372 386512 246424
rect 386564 246412 386570 246424
rect 386564 246384 393314 246412
rect 386564 246372 386570 246384
rect 140774 246304 140780 246356
rect 140832 246344 140838 246356
rect 277486 246344 277492 246356
rect 140832 246316 277492 246344
rect 140832 246304 140838 246316
rect 277486 246304 277492 246316
rect 277544 246304 277550 246356
rect 353478 246304 353484 246356
rect 353536 246344 353542 246356
rect 386414 246344 386420 246356
rect 353536 246316 386420 246344
rect 353536 246304 353542 246316
rect 386414 246304 386420 246316
rect 386472 246304 386478 246356
rect 393286 246344 393314 246384
rect 492674 246344 492680 246356
rect 393286 246316 492680 246344
rect 492674 246304 492680 246316
rect 492732 246304 492738 246356
rect 423030 245556 423036 245608
rect 423088 245596 423094 245608
rect 580166 245596 580172 245608
rect 423088 245568 580172 245596
rect 423088 245556 423094 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 143626 244876 143632 244928
rect 143684 244916 143690 244928
rect 278958 244916 278964 244928
rect 143684 244888 278964 244916
rect 143684 244876 143690 244888
rect 278958 244876 278964 244888
rect 279016 244876 279022 244928
rect 151814 243516 151820 243568
rect 151872 243556 151878 243568
rect 281626 243556 281632 243568
rect 151872 243528 281632 243556
rect 151872 243516 151878 243528
rect 281626 243516 281632 243528
rect 281684 243516 281690 243568
rect 387886 243516 387892 243568
rect 387944 243556 387950 243568
rect 496814 243556 496820 243568
rect 387944 243528 496820 243556
rect 387944 243516 387950 243528
rect 496814 243516 496820 243528
rect 496872 243516 496878 243568
rect 154574 242156 154580 242208
rect 154632 242196 154638 242208
rect 283098 242196 283104 242208
rect 154632 242168 283104 242196
rect 154632 242156 154638 242168
rect 283098 242156 283104 242168
rect 283156 242156 283162 242208
rect 389266 242156 389272 242208
rect 389324 242196 389330 242208
rect 499574 242196 499580 242208
rect 389324 242168 499580 242196
rect 389324 242156 389330 242168
rect 499574 242156 499580 242168
rect 499632 242156 499638 242208
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 232590 241448 232596 241460
rect 3292 241420 232596 241448
rect 3292 241408 3298 241420
rect 232590 241408 232596 241420
rect 232648 241408 232654 241460
rect 230474 240728 230480 240780
rect 230532 240768 230538 240780
rect 305270 240768 305276 240780
rect 230532 240740 305276 240768
rect 230532 240728 230538 240740
rect 305270 240728 305276 240740
rect 305328 240728 305334 240780
rect 390646 240728 390652 240780
rect 390704 240768 390710 240780
rect 503714 240768 503720 240780
rect 390704 240740 503720 240768
rect 390704 240728 390710 240740
rect 503714 240728 503720 240740
rect 503772 240728 503778 240780
rect 158714 239368 158720 239420
rect 158772 239408 158778 239420
rect 283006 239408 283012 239420
rect 158772 239380 283012 239408
rect 158772 239368 158778 239380
rect 283006 239368 283012 239380
rect 283064 239368 283070 239420
rect 392026 239368 392032 239420
rect 392084 239408 392090 239420
rect 510614 239408 510620 239420
rect 392084 239380 510620 239408
rect 392084 239368 392090 239380
rect 510614 239368 510620 239380
rect 510672 239368 510678 239420
rect 166994 238008 167000 238060
rect 167052 238048 167058 238060
rect 285766 238048 285772 238060
rect 167052 238020 285772 238048
rect 167052 238008 167058 238020
rect 285766 238008 285772 238020
rect 285824 238008 285830 238060
rect 394786 238008 394792 238060
rect 394844 238048 394850 238060
rect 517514 238048 517520 238060
rect 394844 238020 517520 238048
rect 394844 238008 394850 238020
rect 517514 238008 517520 238020
rect 517572 238008 517578 238060
rect 180794 236648 180800 236700
rect 180852 236688 180858 236700
rect 289998 236688 290004 236700
rect 180852 236660 290004 236688
rect 180852 236648 180858 236660
rect 289998 236648 290004 236660
rect 290056 236648 290062 236700
rect 396258 236648 396264 236700
rect 396316 236688 396322 236700
rect 521654 236688 521660 236700
rect 396316 236660 521660 236688
rect 396316 236648 396322 236660
rect 521654 236648 521660 236660
rect 521712 236648 521718 236700
rect 187694 235220 187700 235272
rect 187752 235260 187758 235272
rect 292666 235260 292672 235272
rect 187752 235232 292672 235260
rect 187752 235220 187758 235232
rect 292666 235220 292672 235232
rect 292724 235220 292730 235272
rect 396166 235220 396172 235272
rect 396224 235260 396230 235272
rect 524414 235260 524420 235272
rect 396224 235232 524420 235260
rect 396224 235220 396230 235232
rect 524414 235220 524420 235232
rect 524472 235220 524478 235272
rect 191834 233860 191840 233912
rect 191892 233900 191898 233912
rect 294046 233900 294052 233912
rect 191892 233872 294052 233900
rect 191892 233860 191898 233872
rect 294046 233860 294052 233872
rect 294104 233860 294110 233912
rect 397454 233860 397460 233912
rect 397512 233900 397518 233912
rect 528554 233900 528560 233912
rect 397512 233872 528560 233900
rect 397512 233860 397518 233872
rect 528554 233860 528560 233872
rect 528612 233860 528618 233912
rect 429838 233180 429844 233232
rect 429896 233220 429902 233232
rect 579614 233220 579620 233232
rect 429896 233192 579620 233220
rect 429896 233180 429902 233192
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 131114 232500 131120 232552
rect 131172 232540 131178 232552
rect 274726 232540 274732 232552
rect 131172 232512 274732 232540
rect 131172 232500 131178 232512
rect 274726 232500 274732 232512
rect 274784 232500 274790 232552
rect 201586 231072 201592 231124
rect 201644 231112 201650 231124
rect 296806 231112 296812 231124
rect 201644 231084 296812 231112
rect 201644 231072 201650 231084
rect 296806 231072 296812 231084
rect 296864 231072 296870 231124
rect 401778 231072 401784 231124
rect 401836 231112 401842 231124
rect 539594 231112 539600 231124
rect 401836 231084 539600 231112
rect 401836 231072 401842 231084
rect 539594 231072 539600 231084
rect 539652 231072 539658 231124
rect 209866 229712 209872 229764
rect 209924 229752 209930 229764
rect 299658 229752 299664 229764
rect 209924 229724 299664 229752
rect 209924 229712 209930 229724
rect 299658 229712 299664 229724
rect 299716 229712 299722 229764
rect 401686 229712 401692 229764
rect 401744 229752 401750 229764
rect 542354 229752 542360 229764
rect 401744 229724 542360 229752
rect 401744 229712 401750 229724
rect 542354 229712 542360 229724
rect 542412 229712 542418 229764
rect 212534 228352 212540 228404
rect 212592 228392 212598 228404
rect 299566 228392 299572 228404
rect 212592 228364 299572 228392
rect 212592 228352 212598 228364
rect 299566 228352 299572 228364
rect 299624 228352 299630 228404
rect 405826 228352 405832 228404
rect 405884 228392 405890 228404
rect 553394 228392 553400 228404
rect 405884 228364 553400 228392
rect 405884 228352 405890 228364
rect 553394 228352 553400 228364
rect 553452 228352 553458 228404
rect 219434 226992 219440 227044
rect 219492 227032 219498 227044
rect 302418 227032 302424 227044
rect 219492 227004 302424 227032
rect 219492 226992 219498 227004
rect 302418 226992 302424 227004
rect 302476 226992 302482 227044
rect 407206 226992 407212 227044
rect 407264 227032 407270 227044
rect 560294 227032 560300 227044
rect 407264 227004 560300 227032
rect 407264 226992 407270 227004
rect 560294 226992 560300 227004
rect 560352 226992 560358 227044
rect 142154 225564 142160 225616
rect 142212 225604 142218 225616
rect 278866 225604 278872 225616
rect 142212 225576 278872 225604
rect 142212 225564 142218 225576
rect 278866 225564 278872 225576
rect 278924 225564 278930 225616
rect 409966 225564 409972 225616
rect 410024 225604 410030 225616
rect 567194 225604 567200 225616
rect 410024 225576 567200 225604
rect 410024 225564 410030 225576
rect 567194 225564 567200 225576
rect 567252 225564 567258 225616
rect 96614 224204 96620 224256
rect 96672 224244 96678 224256
rect 265158 224244 265164 224256
rect 96672 224216 265164 224244
rect 96672 224204 96678 224216
rect 265158 224204 265164 224216
rect 265216 224204 265222 224256
rect 411346 224204 411352 224256
rect 411404 224244 411410 224256
rect 574094 224244 574100 224256
rect 411404 224216 574100 224244
rect 411404 224204 411410 224216
rect 574094 224204 574100 224216
rect 574152 224204 574158 224256
rect 100754 222844 100760 222896
rect 100812 222884 100818 222896
rect 265066 222884 265072 222896
rect 100812 222856 265072 222884
rect 100812 222844 100818 222856
rect 265066 222844 265072 222856
rect 265124 222844 265130 222896
rect 403618 222844 403624 222896
rect 403676 222884 403682 222896
rect 540974 222884 540980 222896
rect 403676 222856 540980 222884
rect 403676 222844 403682 222856
rect 540974 222844 540980 222856
rect 541032 222844 541038 222896
rect 33134 221416 33140 221468
rect 33192 221456 33198 221468
rect 244458 221456 244464 221468
rect 33192 221428 244464 221456
rect 33192 221416 33198 221428
rect 244458 221416 244464 221428
rect 244516 221416 244522 221468
rect 44174 220056 44180 220108
rect 44232 220096 44238 220108
rect 248598 220096 248604 220108
rect 44232 220068 248604 220096
rect 44232 220056 44238 220068
rect 248598 220056 248604 220068
rect 248656 220056 248662 220108
rect 436738 219376 436744 219428
rect 436796 219416 436802 219428
rect 580166 219416 580172 219428
rect 436796 219388 580172 219416
rect 436796 219376 436802 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 48314 218696 48320 218748
rect 48372 218736 48378 218748
rect 249978 218736 249984 218748
rect 48372 218708 249984 218736
rect 48372 218696 48378 218708
rect 249978 218696 249984 218708
rect 250036 218696 250042 218748
rect 52454 217268 52460 217320
rect 52512 217308 52518 217320
rect 249886 217308 249892 217320
rect 52512 217280 249892 217308
rect 52512 217268 52518 217280
rect 249886 217268 249892 217280
rect 249944 217268 249950 217320
rect 59354 215908 59360 215960
rect 59412 215948 59418 215960
rect 251818 215948 251824 215960
rect 59412 215920 251824 215948
rect 59412 215908 59418 215920
rect 251818 215908 251824 215920
rect 251876 215908 251882 215960
rect 2774 214956 2780 215008
rect 2832 214996 2838 215008
rect 4890 214996 4896 215008
rect 2832 214968 4896 214996
rect 2832 214956 2838 214968
rect 4890 214956 4896 214968
rect 4948 214956 4954 215008
rect 66254 214548 66260 214600
rect 66312 214588 66318 214600
rect 255498 214588 255504 214600
rect 66312 214560 255504 214588
rect 66312 214548 66318 214560
rect 255498 214548 255504 214560
rect 255556 214548 255562 214600
rect 18598 213188 18604 213240
rect 18656 213228 18662 213240
rect 238938 213228 238944 213240
rect 18656 213200 238944 213228
rect 18656 213188 18662 213200
rect 238938 213188 238944 213200
rect 238996 213188 239002 213240
rect 84194 211760 84200 211812
rect 84252 211800 84258 211812
rect 261018 211800 261024 211812
rect 84252 211772 261024 211800
rect 84252 211760 84258 211772
rect 261018 211760 261024 211772
rect 261076 211760 261082 211812
rect 86954 210400 86960 210452
rect 87012 210440 87018 210452
rect 260926 210440 260932 210452
rect 87012 210412 260932 210440
rect 87012 210400 87018 210412
rect 260926 210400 260932 210412
rect 260984 210400 260990 210452
rect 102134 209040 102140 209092
rect 102192 209080 102198 209092
rect 266538 209080 266544 209092
rect 102192 209052 266544 209080
rect 102192 209040 102198 209052
rect 266538 209040 266544 209052
rect 266596 209040 266602 209092
rect 104894 207612 104900 207664
rect 104952 207652 104958 207664
rect 266446 207652 266452 207664
rect 104952 207624 266452 207652
rect 104952 207612 104958 207624
rect 266446 207612 266452 207624
rect 266504 207612 266510 207664
rect 479518 206932 479524 206984
rect 479576 206972 479582 206984
rect 580166 206972 580172 206984
rect 479576 206944 580172 206972
rect 479576 206932 479582 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 27614 206252 27620 206304
rect 27672 206292 27678 206304
rect 242986 206292 242992 206304
rect 27672 206264 242992 206292
rect 27672 206252 27678 206264
rect 242986 206252 242992 206264
rect 243044 206252 243050 206304
rect 30374 204892 30380 204944
rect 30432 204932 30438 204944
rect 244366 204932 244372 204944
rect 30432 204904 244372 204932
rect 30432 204892 30438 204904
rect 244366 204892 244372 204904
rect 244424 204892 244430 204944
rect 13170 203532 13176 203584
rect 13228 203572 13234 203584
rect 237558 203572 237564 203584
rect 13228 203544 237564 203572
rect 13228 203532 13234 203544
rect 237558 203532 237564 203544
rect 237616 203532 237622 203584
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 18690 202824 18696 202836
rect 3384 202796 18696 202824
rect 3384 202784 3390 202796
rect 18690 202784 18696 202796
rect 18748 202784 18754 202836
rect 56594 202104 56600 202156
rect 56652 202144 56658 202156
rect 252646 202144 252652 202156
rect 56652 202116 252652 202144
rect 56652 202104 56658 202116
rect 252646 202104 252652 202116
rect 252704 202104 252710 202156
rect 63494 200744 63500 200796
rect 63552 200784 63558 200796
rect 254210 200784 254216 200796
rect 63552 200756 254216 200784
rect 63552 200744 63558 200756
rect 254210 200744 254216 200756
rect 254268 200744 254274 200796
rect 67634 199384 67640 199436
rect 67692 199424 67698 199436
rect 255406 199424 255412 199436
rect 67692 199396 255412 199424
rect 67692 199384 67698 199396
rect 255406 199384 255412 199396
rect 255464 199384 255470 199436
rect 70394 197956 70400 198008
rect 70452 197996 70458 198008
rect 256878 197996 256884 198008
rect 70452 197968 256884 197996
rect 70452 197956 70458 197968
rect 256878 197956 256884 197968
rect 256936 197956 256942 198008
rect 77294 196596 77300 196648
rect 77352 196636 77358 196648
rect 258258 196636 258264 196648
rect 77352 196608 258264 196636
rect 77352 196596 77358 196608
rect 258258 196596 258264 196608
rect 258316 196596 258322 196648
rect 88334 195236 88340 195288
rect 88392 195276 88398 195288
rect 262398 195276 262404 195288
rect 88392 195248 262404 195276
rect 88392 195236 88398 195248
rect 262398 195236 262404 195248
rect 262456 195236 262462 195288
rect 92474 193808 92480 193860
rect 92532 193848 92538 193860
rect 262306 193848 262312 193860
rect 92532 193820 262312 193848
rect 92532 193808 92538 193820
rect 262306 193808 262312 193820
rect 262364 193808 262370 193860
rect 428458 193128 428464 193180
rect 428516 193168 428522 193180
rect 580166 193168 580172 193180
rect 428516 193140 580172 193168
rect 428516 193128 428522 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 95234 192448 95240 192500
rect 95292 192488 95298 192500
rect 263778 192488 263784 192500
rect 95292 192460 263784 192488
rect 95292 192448 95298 192460
rect 263778 192448 263784 192460
rect 263836 192448 263842 192500
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 11790 189020 11796 189032
rect 3200 188992 11796 189020
rect 3200 188980 3206 188992
rect 11790 188980 11796 188992
rect 11848 188980 11854 189032
rect 263778 180072 263784 180124
rect 263836 180112 263842 180124
rect 316310 180112 316316 180124
rect 263836 180084 316316 180112
rect 263836 180072 263842 180084
rect 316310 180072 316316 180084
rect 316368 180072 316374 180124
rect 435358 179324 435364 179376
rect 435416 179364 435422 179376
rect 580166 179364 580172 179376
rect 435416 179336 580172 179364
rect 435416 179324 435422 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 421558 166948 421564 167000
rect 421616 166988 421622 167000
rect 580166 166988 580172 167000
rect 421616 166960 580172 166988
rect 421616 166948 421622 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 229738 164200 229744 164212
rect 3384 164172 229744 164200
rect 3384 164160 3390 164172
rect 229738 164160 229744 164172
rect 229796 164160 229802 164212
rect 427078 153144 427084 153196
rect 427136 153184 427142 153196
rect 580166 153184 580172 153196
rect 427136 153156 580172 153184
rect 427136 153144 427142 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 21358 150396 21364 150408
rect 3384 150368 21364 150396
rect 3384 150356 3390 150368
rect 21358 150356 21364 150368
rect 21416 150356 21422 150408
rect 424318 139340 424324 139392
rect 424376 139380 424382 139392
rect 580166 139380 580172 139392
rect 424376 139352 580172 139380
rect 424376 139340 424382 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 420178 126896 420184 126948
rect 420236 126936 420242 126948
rect 579614 126936 579620 126948
rect 420236 126908 579620 126936
rect 420236 126896 420242 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 438118 113092 438124 113144
rect 438176 113132 438182 113144
rect 580166 113132 580172 113144
rect 438176 113104 580172 113132
rect 438176 113092 438182 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 432598 100648 432604 100700
rect 432656 100688 432662 100700
rect 579706 100688 579712 100700
rect 432656 100660 579712 100688
rect 432656 100648 432662 100660
rect 579706 100648 579712 100660
rect 579764 100648 579770 100700
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 22738 97968 22744 97980
rect 3568 97940 22744 97968
rect 3568 97928 3574 97940
rect 22738 97928 22744 97940
rect 22796 97928 22802 97980
rect 418798 86912 418804 86964
rect 418856 86952 418862 86964
rect 579982 86952 579988 86964
rect 418856 86924 579988 86952
rect 418856 86912 418862 86924
rect 579982 86912 579988 86924
rect 580040 86912 580046 86964
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 13078 85524 13084 85536
rect 3568 85496 13084 85524
rect 3568 85484 3574 85496
rect 13078 85484 13084 85496
rect 13136 85484 13142 85536
rect 425698 73108 425704 73160
rect 425756 73148 425762 73160
rect 580166 73148 580172 73160
rect 425756 73120 580172 73148
rect 425756 73108 425762 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 44266 72428 44272 72480
rect 44324 72468 44330 72480
rect 248506 72468 248512 72480
rect 44324 72440 248512 72468
rect 44324 72428 44330 72440
rect 248506 72428 248512 72440
rect 248564 72428 248570 72480
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 7558 71652 7564 71664
rect 3568 71624 7564 71652
rect 3568 71612 3574 71624
rect 7558 71612 7564 71624
rect 7616 71612 7622 71664
rect 155954 71000 155960 71052
rect 156012 71040 156018 71052
rect 282914 71040 282920 71052
rect 156012 71012 282920 71040
rect 156012 71000 156018 71012
rect 282914 71000 282920 71012
rect 282972 71000 282978 71052
rect 52546 64132 52552 64184
rect 52604 64172 52610 64184
rect 251266 64172 251272 64184
rect 52604 64144 251272 64172
rect 52604 64132 52610 64144
rect 251266 64132 251272 64144
rect 251324 64132 251330 64184
rect 69106 61344 69112 61396
rect 69164 61384 69170 61396
rect 255314 61384 255320 61396
rect 69164 61356 255320 61384
rect 69164 61344 69170 61356
rect 255314 61344 255320 61356
rect 255372 61344 255378 61396
rect 431218 60664 431224 60716
rect 431276 60704 431282 60716
rect 579798 60704 579804 60716
rect 431276 60676 579804 60704
rect 431276 60664 431282 60676
rect 579798 60664 579804 60676
rect 579856 60664 579862 60716
rect 97994 59984 98000 60036
rect 98052 60024 98058 60036
rect 265250 60024 265256 60036
rect 98052 59996 265256 60024
rect 98052 59984 98058 59996
rect 265250 59984 265256 59996
rect 265308 59984 265314 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 10410 59344 10416 59356
rect 3108 59316 10416 59344
rect 3108 59304 3114 59316
rect 10410 59304 10416 59316
rect 10468 59304 10474 59356
rect 85666 55836 85672 55888
rect 85724 55876 85730 55888
rect 260834 55876 260840 55888
rect 85724 55848 260840 55876
rect 85724 55836 85730 55848
rect 260834 55836 260840 55848
rect 260892 55836 260898 55888
rect 160186 54476 160192 54528
rect 160244 54516 160250 54528
rect 284386 54516 284392 54528
rect 160244 54488 284392 54516
rect 160244 54476 160250 54488
rect 284386 54476 284392 54488
rect 284444 54476 284450 54528
rect 151906 53048 151912 53100
rect 151964 53088 151970 53100
rect 281534 53088 281540 53100
rect 151964 53060 281540 53088
rect 151964 53048 151970 53060
rect 281534 53048 281540 53060
rect 281592 53048 281598 53100
rect 138014 51688 138020 51740
rect 138072 51728 138078 51740
rect 277670 51728 277676 51740
rect 138072 51700 277676 51728
rect 138072 51688 138078 51700
rect 277670 51688 277676 51700
rect 277728 51688 277734 51740
rect 347958 51688 347964 51740
rect 348016 51728 348022 51740
rect 365806 51728 365812 51740
rect 348016 51700 365812 51728
rect 348016 51688 348022 51700
rect 365806 51688 365812 51700
rect 365864 51688 365870 51740
rect 149054 50328 149060 50380
rect 149112 50368 149118 50380
rect 280154 50368 280160 50380
rect 149112 50340 280160 50368
rect 149112 50328 149118 50340
rect 280154 50328 280160 50340
rect 280212 50328 280218 50380
rect 2774 48968 2780 49020
rect 2832 49008 2838 49020
rect 234614 49008 234620 49020
rect 2832 48980 234620 49008
rect 2832 48968 2838 48980
rect 234614 48968 234620 48980
rect 234672 48968 234678 49020
rect 251266 48968 251272 49020
rect 251324 49008 251330 49020
rect 312078 49008 312084 49020
rect 251324 48980 312084 49008
rect 251324 48968 251330 48980
rect 312078 48968 312084 48980
rect 312136 48968 312142 49020
rect 244366 47540 244372 47592
rect 244424 47580 244430 47592
rect 310698 47580 310704 47592
rect 244424 47552 310704 47580
rect 244424 47540 244430 47552
rect 310698 47540 310704 47552
rect 310756 47540 310762 47592
rect 353386 47540 353392 47592
rect 353444 47580 353450 47592
rect 385126 47580 385132 47592
rect 353444 47552 385132 47580
rect 353444 47540 353450 47552
rect 385126 47540 385132 47552
rect 385184 47540 385190 47592
rect 417418 46860 417424 46912
rect 417476 46900 417482 46912
rect 580166 46900 580172 46912
rect 417476 46872 580172 46900
rect 417476 46860 417482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 241698 46180 241704 46232
rect 241756 46220 241762 46232
rect 309318 46220 309324 46232
rect 241756 46192 309324 46220
rect 241756 46180 241762 46192
rect 309318 46180 309324 46192
rect 309376 46180 309382 46232
rect 237558 44820 237564 44872
rect 237616 44860 237622 44872
rect 307846 44860 307852 44872
rect 237616 44832 307852 44860
rect 237616 44820 237622 44832
rect 307846 44820 307852 44832
rect 307904 44820 307910 44872
rect 135346 43392 135352 43444
rect 135404 43432 135410 43444
rect 276014 43432 276020 43444
rect 135404 43404 276020 43432
rect 135404 43392 135410 43404
rect 276014 43392 276020 43404
rect 276072 43392 276078 43444
rect 194594 42032 194600 42084
rect 194652 42072 194658 42084
rect 294230 42072 294236 42084
rect 194652 42044 294236 42072
rect 194652 42032 194658 42044
rect 294230 42032 294236 42044
rect 294288 42032 294294 42084
rect 398834 42032 398840 42084
rect 398892 42072 398898 42084
rect 531406 42072 531412 42084
rect 398892 42044 531412 42072
rect 398892 42032 398898 42044
rect 531406 42032 531412 42044
rect 531464 42032 531470 42084
rect 185026 40672 185032 40724
rect 185084 40712 185090 40724
rect 291470 40712 291476 40724
rect 185084 40684 291476 40712
rect 185084 40672 185090 40684
rect 291470 40672 291476 40684
rect 291528 40672 291534 40724
rect 198734 39312 198740 39364
rect 198792 39352 198798 39364
rect 295334 39352 295340 39364
rect 198792 39324 295340 39352
rect 198792 39312 198798 39324
rect 295334 39312 295340 39324
rect 295392 39312 295398 39364
rect 169754 37884 169760 37936
rect 169812 37924 169818 37936
rect 287330 37924 287336 37936
rect 169812 37896 287336 37924
rect 169812 37884 169818 37896
rect 287330 37884 287336 37896
rect 287388 37884 287394 37936
rect 162854 36524 162860 36576
rect 162912 36564 162918 36576
rect 284570 36564 284576 36576
rect 162912 36536 284576 36564
rect 162912 36524 162918 36536
rect 284570 36524 284576 36536
rect 284628 36524 284634 36576
rect 411254 36524 411260 36576
rect 411312 36564 411318 36576
rect 571334 36564 571340 36576
rect 411312 36536 571340 36564
rect 411312 36524 411318 36536
rect 571334 36524 571340 36536
rect 571392 36524 571398 36576
rect 126974 35164 126980 35216
rect 127032 35204 127038 35216
rect 273346 35204 273352 35216
rect 127032 35176 273352 35204
rect 127032 35164 127038 35176
rect 273346 35164 273352 35176
rect 273404 35164 273410 35216
rect 282914 35164 282920 35216
rect 282972 35204 282978 35216
rect 307018 35204 307024 35216
rect 282972 35176 307024 35204
rect 282972 35164 282978 35176
rect 307018 35164 307024 35176
rect 307076 35164 307082 35216
rect 73154 33736 73160 33788
rect 73212 33776 73218 33788
rect 256786 33776 256792 33788
rect 73212 33748 256792 33776
rect 73212 33736 73218 33748
rect 256786 33736 256792 33748
rect 256844 33736 256850 33788
rect 264974 33736 264980 33788
rect 265032 33776 265038 33788
rect 316218 33776 316224 33788
rect 265032 33748 316224 33776
rect 265032 33736 265038 33748
rect 316218 33736 316224 33748
rect 316276 33736 316282 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 8938 33096 8944 33108
rect 3568 33068 8944 33096
rect 3568 33056 3574 33068
rect 8938 33056 8944 33068
rect 8996 33056 9002 33108
rect 55214 32376 55220 32428
rect 55272 32416 55278 32428
rect 251174 32416 251180 32428
rect 55272 32388 251180 32416
rect 55272 32376 55278 32388
rect 251174 32376 251180 32388
rect 251232 32376 251238 32428
rect 258258 32376 258264 32428
rect 258316 32416 258322 32428
rect 314746 32416 314752 32428
rect 258316 32388 314752 32416
rect 258316 32376 258322 32388
rect 314746 32376 314752 32388
rect 314804 32376 314810 32428
rect 357526 32376 357532 32428
rect 357584 32416 357590 32428
rect 397454 32416 397460 32428
rect 357584 32388 397460 32416
rect 357584 32376 357590 32388
rect 397454 32376 397460 32388
rect 397512 32376 397518 32428
rect 400214 32376 400220 32428
rect 400272 32416 400278 32428
rect 535454 32416 535460 32428
rect 400272 32388 535460 32416
rect 400272 32376 400278 32388
rect 535454 32376 535460 32388
rect 535512 32376 535518 32428
rect 49694 31016 49700 31068
rect 49752 31056 49758 31068
rect 249794 31056 249800 31068
rect 49752 31028 249800 31056
rect 49752 31016 49758 31028
rect 249794 31016 249800 31028
rect 249852 31016 249858 31068
rect 251174 31016 251180 31068
rect 251232 31056 251238 31068
rect 311986 31056 311992 31068
rect 251232 31028 311992 31056
rect 251232 31016 251238 31028
rect 311986 31016 311992 31028
rect 312044 31016 312050 31068
rect 358906 31016 358912 31068
rect 358964 31056 358970 31068
rect 404446 31056 404452 31068
rect 358964 31028 404452 31056
rect 358964 31016 358970 31028
rect 404446 31016 404452 31028
rect 404504 31016 404510 31068
rect 247218 29656 247224 29708
rect 247276 29696 247282 29708
rect 310606 29696 310612 29708
rect 247276 29668 310612 29696
rect 247276 29656 247282 29668
rect 310606 29656 310612 29668
rect 310664 29656 310670 29708
rect 60826 29588 60832 29640
rect 60884 29628 60890 29640
rect 252738 29628 252744 29640
rect 60884 29600 252744 29628
rect 60884 29588 60890 29600
rect 252738 29588 252744 29600
rect 252796 29588 252802 29640
rect 310698 29588 310704 29640
rect 310756 29628 310762 29640
rect 330110 29628 330116 29640
rect 310756 29600 330116 29628
rect 310756 29588 310762 29600
rect 330110 29588 330116 29600
rect 330168 29588 330174 29640
rect 354766 29588 354772 29640
rect 354824 29628 354830 29640
rect 390738 29628 390744 29640
rect 354824 29600 390744 29628
rect 354824 29588 354830 29600
rect 390738 29588 390744 29600
rect 390796 29588 390802 29640
rect 408494 29588 408500 29640
rect 408552 29628 408558 29640
rect 564526 29628 564532 29640
rect 408552 29600 564532 29628
rect 408552 29588 408558 29600
rect 564526 29588 564532 29600
rect 564584 29588 564590 29640
rect 356146 28364 356152 28416
rect 356204 28404 356210 28416
rect 393406 28404 393412 28416
rect 356204 28376 393412 28404
rect 356204 28364 356210 28376
rect 393406 28364 393412 28376
rect 393464 28364 393470 28416
rect 242986 28228 242992 28280
rect 243044 28268 243050 28280
rect 309226 28268 309232 28280
rect 243044 28240 309232 28268
rect 243044 28228 243050 28240
rect 309226 28228 309232 28240
rect 309284 28228 309290 28280
rect 393314 28228 393320 28280
rect 393372 28268 393378 28280
rect 514846 28268 514852 28280
rect 393372 28240 514852 28268
rect 393372 28228 393378 28240
rect 514846 28228 514852 28240
rect 514904 28228 514910 28280
rect 240318 26868 240324 26920
rect 240376 26908 240382 26920
rect 309410 26908 309416 26920
rect 240376 26880 309416 26908
rect 240376 26868 240382 26880
rect 309410 26868 309416 26880
rect 309468 26868 309474 26920
rect 350626 26868 350632 26920
rect 350684 26908 350690 26920
rect 375558 26908 375564 26920
rect 350684 26880 375564 26908
rect 350684 26868 350690 26880
rect 375558 26868 375564 26880
rect 375616 26868 375622 26920
rect 390554 26868 390560 26920
rect 390612 26908 390618 26920
rect 506566 26908 506572 26920
rect 390612 26880 506572 26908
rect 390612 26868 390618 26880
rect 506566 26868 506572 26880
rect 506624 26868 506630 26920
rect 262306 25576 262312 25628
rect 262364 25616 262370 25628
rect 316126 25616 316132 25628
rect 262364 25588 316132 25616
rect 262364 25576 262370 25588
rect 316126 25576 316132 25588
rect 316184 25576 316190 25628
rect 218054 25508 218060 25560
rect 218112 25548 218118 25560
rect 298738 25548 298744 25560
rect 218112 25520 298744 25548
rect 218112 25508 218118 25520
rect 298738 25508 298744 25520
rect 298796 25508 298802 25560
rect 358078 25508 358084 25560
rect 358136 25548 358142 25560
rect 372798 25548 372804 25560
rect 358136 25520 372804 25548
rect 358136 25508 358142 25520
rect 372798 25508 372804 25520
rect 372856 25508 372862 25560
rect 385034 25508 385040 25560
rect 385092 25548 385098 25560
rect 490006 25548 490012 25560
rect 385092 25520 490012 25548
rect 385092 25508 385098 25520
rect 490006 25508 490012 25520
rect 490064 25508 490070 25560
rect 268010 24148 268016 24200
rect 268068 24188 268074 24200
rect 317598 24188 317604 24200
rect 268068 24160 317604 24188
rect 268068 24148 268074 24160
rect 317598 24148 317604 24160
rect 317656 24148 317662 24200
rect 127066 24080 127072 24132
rect 127124 24120 127130 24132
rect 273530 24120 273536 24132
rect 127124 24092 273536 24120
rect 127124 24080 127130 24092
rect 273530 24080 273536 24092
rect 273588 24080 273594 24132
rect 360378 24080 360384 24132
rect 360436 24120 360442 24132
rect 407206 24120 407212 24132
rect 360436 24092 407212 24120
rect 360436 24080 360442 24092
rect 407206 24080 407212 24092
rect 407264 24080 407270 24132
rect 256786 22788 256792 22840
rect 256844 22828 256850 22840
rect 313366 22828 313372 22840
rect 256844 22800 313372 22828
rect 256844 22788 256850 22800
rect 313366 22788 313372 22800
rect 313424 22788 313430 22840
rect 144914 22720 144920 22772
rect 144972 22760 144978 22772
rect 278774 22760 278780 22772
rect 144972 22732 278780 22760
rect 144972 22720 144978 22732
rect 278774 22720 278780 22732
rect 278832 22720 278838 22772
rect 356054 22720 356060 22772
rect 356112 22760 356118 22772
rect 396166 22760 396172 22772
rect 356112 22732 396172 22760
rect 356112 22720 356118 22732
rect 396166 22720 396172 22732
rect 396224 22720 396230 22772
rect 37274 21360 37280 21412
rect 37332 21400 37338 21412
rect 245746 21400 245752 21412
rect 37332 21372 245752 21400
rect 37332 21360 37338 21372
rect 245746 21360 245752 21372
rect 245804 21360 245810 21412
rect 252554 21360 252560 21412
rect 252612 21400 252618 21412
rect 312170 21400 312176 21412
rect 252612 21372 312176 21400
rect 252612 21360 252618 21372
rect 312170 21360 312176 21372
rect 312228 21360 312234 21412
rect 352098 21360 352104 21412
rect 352156 21400 352162 21412
rect 382458 21400 382464 21412
rect 352156 21372 382464 21400
rect 352156 21360 352162 21372
rect 382458 21360 382464 21372
rect 382516 21360 382522 21412
rect 396074 21360 396080 21412
rect 396132 21400 396138 21412
rect 523034 21400 523040 21412
rect 396132 21372 523040 21400
rect 396132 21360 396138 21372
rect 523034 21360 523040 21372
rect 523092 21360 523098 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 414934 20652 414940 20664
rect 3476 20624 414940 20652
rect 3476 20612 3482 20624
rect 414934 20612 414940 20624
rect 414992 20612 414998 20664
rect 259730 19932 259736 19984
rect 259788 19972 259794 19984
rect 302970 19972 302976 19984
rect 259788 19944 302976 19972
rect 259788 19932 259794 19944
rect 302970 19932 302976 19944
rect 303028 19932 303034 19984
rect 248506 18640 248512 18692
rect 248564 18680 248570 18692
rect 310790 18680 310796 18692
rect 248564 18652 310796 18680
rect 248564 18640 248570 18652
rect 310790 18640 310796 18652
rect 310848 18640 310854 18692
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 238846 18612 238852 18624
rect 13872 18584 238852 18612
rect 13872 18572 13878 18584
rect 238846 18572 238852 18584
rect 238904 18572 238910 18624
rect 238938 18572 238944 18624
rect 238996 18612 239002 18624
rect 301498 18612 301504 18624
rect 238996 18584 301504 18612
rect 238996 18572 239002 18584
rect 301498 18572 301504 18584
rect 301556 18572 301562 18624
rect 307754 18572 307760 18624
rect 307812 18612 307818 18624
rect 330018 18612 330024 18624
rect 307812 18584 330024 18612
rect 307812 18572 307818 18584
rect 330018 18572 330024 18584
rect 330076 18572 330082 18624
rect 347866 18572 347872 18624
rect 347924 18612 347930 18624
rect 368750 18612 368756 18624
rect 347924 18584 368756 18612
rect 347924 18572 347930 18584
rect 368750 18572 368756 18584
rect 368808 18572 368814 18624
rect 370498 18572 370504 18624
rect 370556 18612 370562 18624
rect 412818 18612 412824 18624
rect 370556 18584 412824 18612
rect 370556 18572 370562 18584
rect 412818 18572 412824 18584
rect 412876 18572 412882 18624
rect 234614 17348 234620 17400
rect 234672 17388 234678 17400
rect 306650 17388 306656 17400
rect 234672 17360 306656 17388
rect 234672 17348 234678 17360
rect 306650 17348 306656 17360
rect 306708 17348 306714 17400
rect 360286 17348 360292 17400
rect 360344 17388 360350 17400
rect 405826 17388 405832 17400
rect 360344 17360 405832 17388
rect 360344 17348 360350 17360
rect 405826 17348 405832 17360
rect 405884 17348 405890 17400
rect 255314 17280 255320 17332
rect 255372 17320 255378 17332
rect 313458 17320 313464 17332
rect 255372 17292 313464 17320
rect 255372 17280 255378 17292
rect 313458 17280 313464 17292
rect 313516 17280 313522 17332
rect 306466 17212 306472 17264
rect 306524 17252 306530 17264
rect 328638 17252 328644 17264
rect 306524 17224 328644 17252
rect 306524 17212 306530 17224
rect 328638 17212 328644 17224
rect 328696 17212 328702 17264
rect 346578 17212 346584 17264
rect 346636 17252 346642 17264
rect 360286 17252 360292 17264
rect 346636 17224 360292 17252
rect 346636 17212 346642 17224
rect 360286 17212 360292 17224
rect 360344 17212 360350 17264
rect 405734 17212 405740 17264
rect 405792 17252 405798 17264
rect 556246 17252 556252 17264
rect 405792 17224 556252 17252
rect 405792 17212 405798 17224
rect 556246 17212 556252 17224
rect 556304 17212 556310 17264
rect 260650 15920 260656 15972
rect 260708 15960 260714 15972
rect 291838 15960 291844 15972
rect 260708 15932 291844 15960
rect 260708 15920 260714 15932
rect 291838 15920 291844 15932
rect 291896 15920 291902 15972
rect 116394 15852 116400 15904
rect 116452 15892 116458 15904
rect 270678 15892 270684 15904
rect 116452 15864 270684 15892
rect 116452 15852 116458 15864
rect 270678 15852 270684 15864
rect 270736 15852 270742 15904
rect 279050 15852 279056 15904
rect 279108 15892 279114 15904
rect 319438 15892 319444 15904
rect 279108 15864 319444 15892
rect 279108 15852 279114 15864
rect 319438 15852 319444 15864
rect 319496 15852 319502 15904
rect 358814 15852 358820 15904
rect 358872 15892 358878 15904
rect 402514 15892 402520 15904
rect 358872 15864 402520 15892
rect 358872 15852 358878 15864
rect 402514 15852 402520 15864
rect 402572 15852 402578 15904
rect 404354 15852 404360 15904
rect 404412 15892 404418 15904
rect 550266 15892 550272 15904
rect 404412 15864 550272 15892
rect 404412 15852 404418 15864
rect 550266 15852 550272 15864
rect 550324 15852 550330 15904
rect 112346 14764 112352 14816
rect 112404 14804 112410 14816
rect 269298 14804 269304 14816
rect 112404 14776 269304 14804
rect 112404 14764 112410 14776
rect 269298 14764 269304 14776
rect 269356 14764 269362 14816
rect 109034 14696 109040 14748
rect 109092 14736 109098 14748
rect 267918 14736 267924 14748
rect 109092 14708 267924 14736
rect 109092 14696 109098 14708
rect 267918 14696 267924 14708
rect 267976 14696 267982 14748
rect 93854 14628 93860 14680
rect 93912 14668 93918 14680
rect 263686 14668 263692 14680
rect 93912 14640 263692 14668
rect 93912 14628 93918 14640
rect 263686 14628 263692 14640
rect 263744 14628 263750 14680
rect 91554 14560 91560 14612
rect 91612 14600 91618 14612
rect 262214 14600 262220 14612
rect 91612 14572 262220 14600
rect 91612 14560 91618 14572
rect 262214 14560 262220 14572
rect 262272 14560 262278 14612
rect 80882 14492 80888 14544
rect 80940 14532 80946 14544
rect 259638 14532 259644 14544
rect 80940 14504 259644 14532
rect 80940 14492 80946 14504
rect 259638 14492 259644 14504
rect 259696 14492 259702 14544
rect 313826 14492 313832 14544
rect 313884 14532 313890 14544
rect 331490 14532 331496 14544
rect 313884 14504 331496 14532
rect 313884 14492 313890 14504
rect 331490 14492 331496 14504
rect 331548 14492 331554 14544
rect 77386 14424 77392 14476
rect 77444 14464 77450 14476
rect 258166 14464 258172 14476
rect 77444 14436 258172 14464
rect 77444 14424 77450 14436
rect 258166 14424 258172 14436
rect 258224 14424 258230 14476
rect 268102 14424 268108 14476
rect 268160 14464 268166 14476
rect 313918 14464 313924 14476
rect 268160 14436 313924 14464
rect 268160 14424 268166 14436
rect 313918 14424 313924 14436
rect 313976 14424 313982 14476
rect 352006 14424 352012 14476
rect 352064 14464 352070 14476
rect 381170 14464 381176 14476
rect 352064 14436 381176 14464
rect 352064 14424 352070 14436
rect 381170 14424 381176 14436
rect 381228 14424 381234 14476
rect 383654 14424 383660 14476
rect 383712 14464 383718 14476
rect 482370 14464 482376 14476
rect 383712 14436 482376 14464
rect 383712 14424 383718 14436
rect 482370 14424 482376 14436
rect 482428 14424 482434 14476
rect 118786 13336 118792 13388
rect 118844 13376 118850 13388
rect 270770 13376 270776 13388
rect 118844 13348 270776 13376
rect 118844 13336 118850 13348
rect 270770 13336 270776 13348
rect 270828 13336 270834 13388
rect 114738 13268 114744 13320
rect 114796 13308 114802 13320
rect 270586 13308 270592 13320
rect 114796 13280 270592 13308
rect 114796 13268 114802 13280
rect 270586 13268 270592 13280
rect 270644 13268 270650 13320
rect 111610 13200 111616 13252
rect 111668 13240 111674 13252
rect 269206 13240 269212 13252
rect 111668 13212 269212 13240
rect 111668 13200 111674 13212
rect 269206 13200 269212 13212
rect 269264 13200 269270 13252
rect 108114 13132 108120 13184
rect 108172 13172 108178 13184
rect 267826 13172 267832 13184
rect 108172 13144 267832 13172
rect 108172 13132 108178 13144
rect 267826 13132 267832 13144
rect 267884 13132 267890 13184
rect 363046 13132 363052 13184
rect 363104 13172 363110 13184
rect 415486 13172 415492 13184
rect 363104 13144 415492 13172
rect 363104 13132 363110 13144
rect 415486 13132 415492 13144
rect 415544 13132 415550 13184
rect 93946 13064 93952 13116
rect 94004 13104 94010 13116
rect 263594 13104 263600 13116
rect 94004 13076 263600 13104
rect 94004 13064 94010 13076
rect 263594 13064 263600 13076
rect 263652 13064 263658 13116
rect 270770 13064 270776 13116
rect 270828 13104 270834 13116
rect 317506 13104 317512 13116
rect 270828 13076 317512 13104
rect 270828 13064 270834 13076
rect 317506 13064 317512 13076
rect 317564 13064 317570 13116
rect 350534 13064 350540 13116
rect 350592 13104 350598 13116
rect 377306 13104 377312 13116
rect 350592 13076 377312 13104
rect 350592 13064 350598 13076
rect 377306 13064 377312 13076
rect 377364 13064 377370 13116
rect 407114 13064 407120 13116
rect 407172 13104 407178 13116
rect 559282 13104 559288 13116
rect 407172 13076 559288 13104
rect 407172 13064 407178 13076
rect 559282 13064 559288 13076
rect 559340 13064 559346 13116
rect 126974 11772 126980 11824
rect 127032 11812 127038 11824
rect 128170 11812 128176 11824
rect 127032 11784 128176 11812
rect 127032 11772 127038 11784
rect 128170 11772 128176 11784
rect 128228 11772 128234 11824
rect 160094 11772 160100 11824
rect 160152 11812 160158 11824
rect 161290 11812 161296 11824
rect 160152 11784 161296 11812
rect 160152 11772 160158 11784
rect 161290 11772 161296 11784
rect 161348 11772 161354 11824
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 216858 11772 216864 11824
rect 216916 11812 216922 11824
rect 300854 11812 300860 11824
rect 216916 11784 300860 11812
rect 216916 11772 216922 11784
rect 300854 11772 300860 11784
rect 300912 11772 300918 11824
rect 349338 11772 349344 11824
rect 349396 11812 349402 11824
rect 374270 11812 374276 11824
rect 349396 11784 374276 11812
rect 349396 11772 349402 11784
rect 374270 11772 374276 11784
rect 374328 11772 374334 11824
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 237466 11744 237472 11756
rect 8812 11716 237472 11744
rect 8812 11704 8818 11716
rect 237466 11704 237472 11716
rect 237524 11704 237530 11756
rect 271966 11704 271972 11756
rect 272024 11744 272030 11756
rect 318886 11744 318892 11756
rect 272024 11716 318892 11744
rect 272024 11704 272030 11716
rect 318886 11704 318892 11716
rect 318944 11704 318950 11756
rect 373258 11704 373264 11756
rect 373316 11744 373322 11756
rect 414290 11744 414296 11756
rect 373316 11716 414296 11744
rect 373316 11704 373322 11716
rect 414290 11704 414296 11716
rect 414348 11704 414354 11756
rect 422938 11704 422944 11756
rect 422996 11744 423002 11756
rect 523126 11744 523132 11756
rect 422996 11716 523132 11744
rect 422996 11704 423002 11716
rect 523126 11704 523132 11716
rect 523184 11704 523190 11756
rect 226334 11636 226340 11688
rect 226392 11676 226398 11688
rect 227530 11676 227536 11688
rect 226392 11648 227536 11676
rect 226392 11636 226398 11648
rect 227530 11636 227536 11648
rect 227588 11636 227594 11688
rect 372706 10820 372712 10872
rect 372764 10860 372770 10872
rect 445754 10860 445760 10872
rect 372764 10832 445760 10860
rect 372764 10820 372770 10832
rect 445754 10820 445760 10832
rect 445812 10820 445818 10872
rect 372614 10752 372620 10804
rect 372672 10792 372678 10804
rect 448606 10792 448612 10804
rect 372672 10764 448612 10792
rect 372672 10752 372678 10764
rect 448606 10752 448612 10764
rect 448664 10752 448670 10804
rect 374178 10684 374184 10736
rect 374236 10724 374242 10736
rect 453298 10724 453304 10736
rect 374236 10696 453304 10724
rect 374236 10684 374242 10696
rect 453298 10684 453304 10696
rect 453356 10684 453362 10736
rect 375466 10616 375472 10668
rect 375524 10656 375530 10668
rect 456886 10656 456892 10668
rect 375524 10628 456892 10656
rect 375524 10616 375530 10628
rect 456886 10616 456892 10628
rect 456944 10616 456950 10668
rect 376754 10548 376760 10600
rect 376812 10588 376818 10600
rect 459922 10588 459928 10600
rect 376812 10560 459928 10588
rect 376812 10548 376818 10560
rect 459922 10548 459928 10560
rect 459980 10548 459986 10600
rect 378318 10480 378324 10532
rect 378376 10520 378382 10532
rect 463970 10520 463976 10532
rect 378376 10492 463976 10520
rect 378376 10480 378382 10492
rect 463970 10480 463976 10492
rect 464028 10480 464034 10532
rect 173894 10412 173900 10464
rect 173952 10452 173958 10464
rect 288526 10452 288532 10464
rect 173952 10424 288532 10452
rect 173952 10412 173958 10424
rect 288526 10412 288532 10424
rect 288584 10412 288590 10464
rect 378226 10412 378232 10464
rect 378284 10452 378290 10464
rect 467466 10452 467472 10464
rect 378284 10424 467472 10452
rect 378284 10412 378290 10424
rect 467466 10412 467472 10424
rect 467524 10412 467530 10464
rect 83274 10344 83280 10396
rect 83332 10384 83338 10396
rect 259454 10384 259460 10396
rect 83332 10356 259460 10384
rect 83332 10344 83338 10356
rect 259454 10344 259460 10356
rect 259512 10344 259518 10396
rect 345106 10344 345112 10396
rect 345164 10384 345170 10396
rect 357526 10384 357532 10396
rect 345164 10356 357532 10384
rect 345164 10344 345170 10356
rect 357526 10344 357532 10356
rect 357584 10344 357590 10396
rect 380986 10344 380992 10396
rect 381044 10384 381050 10396
rect 474090 10384 474096 10396
rect 381044 10356 474096 10384
rect 381044 10344 381050 10356
rect 474090 10344 474096 10356
rect 474148 10344 474154 10396
rect 79226 10276 79232 10328
rect 79284 10316 79290 10328
rect 259546 10316 259552 10328
rect 79284 10288 259552 10316
rect 79284 10276 79290 10288
rect 259546 10276 259552 10288
rect 259604 10276 259610 10328
rect 261754 10276 261760 10328
rect 261812 10316 261818 10328
rect 314838 10316 314844 10328
rect 261812 10288 314844 10316
rect 261812 10276 261818 10288
rect 314838 10276 314844 10288
rect 314896 10276 314902 10328
rect 349246 10276 349252 10328
rect 349304 10316 349310 10328
rect 371510 10316 371516 10328
rect 349304 10288 371516 10316
rect 349304 10276 349310 10288
rect 371510 10276 371516 10288
rect 371568 10276 371574 10328
rect 382366 10276 382372 10328
rect 382424 10316 382430 10328
rect 478138 10316 478144 10328
rect 382424 10288 478144 10316
rect 382424 10276 382430 10288
rect 478138 10276 478144 10288
rect 478196 10276 478202 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 249978 9120 249984 9172
rect 250036 9160 250042 9172
rect 297358 9160 297364 9172
rect 250036 9132 297364 9160
rect 250036 9120 250042 9132
rect 297358 9120 297364 9132
rect 297416 9120 297422 9172
rect 254670 9052 254676 9104
rect 254728 9092 254734 9104
rect 305730 9092 305736 9104
rect 254728 9064 305736 9092
rect 254728 9052 254734 9064
rect 305730 9052 305736 9064
rect 305788 9052 305794 9104
rect 76190 8984 76196 9036
rect 76248 9024 76254 9036
rect 258074 9024 258080 9036
rect 76248 8996 258080 9024
rect 76248 8984 76254 8996
rect 258074 8984 258080 8996
rect 258132 8984 258138 9036
rect 349154 8984 349160 9036
rect 349212 9024 349218 9036
rect 370590 9024 370596 9036
rect 349212 8996 370596 9024
rect 349212 8984 349218 8996
rect 370590 8984 370596 8996
rect 370648 8984 370654 9036
rect 72602 8916 72608 8968
rect 72660 8956 72666 8968
rect 256694 8956 256700 8968
rect 72660 8928 256700 8956
rect 72660 8916 72666 8928
rect 256694 8916 256700 8928
rect 256752 8916 256758 8968
rect 317322 8916 317328 8968
rect 317380 8956 317386 8968
rect 332778 8956 332784 8968
rect 317380 8928 332784 8956
rect 317380 8916 317386 8928
rect 332778 8916 332784 8928
rect 332836 8916 332842 8968
rect 353294 8916 353300 8968
rect 353352 8956 353358 8968
rect 383562 8956 383568 8968
rect 353352 8928 383568 8956
rect 353352 8916 353358 8928
rect 383562 8916 383568 8928
rect 383620 8916 383626 8968
rect 387058 8916 387064 8968
rect 387116 8956 387122 8968
rect 398834 8956 398840 8968
rect 387116 8928 398840 8956
rect 387116 8916 387122 8928
rect 398834 8916 398840 8928
rect 398892 8916 398898 8968
rect 412726 8916 412732 8968
rect 412784 8956 412790 8968
rect 577406 8956 577412 8968
rect 412784 8928 577412 8956
rect 412784 8916 412790 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 377398 8236 377404 8288
rect 377456 8276 377462 8288
rect 378870 8276 378876 8288
rect 377456 8248 378876 8276
rect 377456 8236 377462 8248
rect 378870 8236 378876 8248
rect 378928 8236 378934 8288
rect 237006 7624 237012 7676
rect 237064 7664 237070 7676
rect 304258 7664 304264 7676
rect 237064 7636 304264 7664
rect 237064 7624 237070 7636
rect 304258 7624 304264 7636
rect 304316 7624 304322 7676
rect 310238 7624 310244 7676
rect 310296 7664 310302 7676
rect 329926 7664 329932 7676
rect 310296 7636 329932 7664
rect 310296 7624 310302 7636
rect 329926 7624 329932 7636
rect 329984 7624 329990 7676
rect 347774 7624 347780 7676
rect 347832 7664 347838 7676
rect 367002 7664 367008 7676
rect 347832 7636 367008 7664
rect 347832 7624 347838 7636
rect 367002 7624 367008 7636
rect 367060 7624 367066 7676
rect 176746 7556 176752 7608
rect 176804 7596 176810 7608
rect 288618 7596 288624 7608
rect 176804 7568 288624 7596
rect 176804 7556 176810 7568
rect 288618 7556 288624 7568
rect 288676 7556 288682 7608
rect 290182 7556 290188 7608
rect 290240 7596 290246 7608
rect 315298 7596 315304 7608
rect 290240 7568 315304 7596
rect 290240 7556 290246 7568
rect 315298 7556 315304 7568
rect 315356 7556 315362 7608
rect 351914 7556 351920 7608
rect 351972 7596 351978 7608
rect 379974 7596 379980 7608
rect 351972 7568 379980 7596
rect 351972 7556 351978 7568
rect 379974 7556 379980 7568
rect 380032 7556 380038 7608
rect 380894 7556 380900 7608
rect 380952 7596 380958 7608
rect 476942 7596 476948 7608
rect 380952 7568 476948 7596
rect 380952 7556 380958 7568
rect 476942 7556 476948 7568
rect 477000 7556 477006 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 14458 6848 14464 6860
rect 3476 6820 14464 6848
rect 3476 6808 3482 6820
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 367186 6468 367192 6520
rect 367244 6508 367250 6520
rect 430850 6508 430856 6520
rect 367244 6480 430856 6508
rect 367244 6468 367250 6480
rect 430850 6468 430856 6480
rect 430908 6468 430914 6520
rect 368658 6400 368664 6452
rect 368716 6440 368722 6452
rect 434438 6440 434444 6452
rect 368716 6412 434444 6440
rect 368716 6400 368722 6412
rect 434438 6400 434444 6412
rect 434496 6400 434502 6452
rect 369946 6332 369952 6384
rect 370004 6372 370010 6384
rect 437934 6372 437940 6384
rect 370004 6344 437940 6372
rect 370004 6332 370010 6344
rect 437934 6332 437940 6344
rect 437992 6332 437998 6384
rect 281902 6264 281908 6316
rect 281960 6304 281966 6316
rect 321738 6304 321744 6316
rect 281960 6276 321744 6304
rect 281960 6264 281966 6276
rect 321738 6264 321744 6276
rect 321796 6264 321802 6316
rect 371326 6264 371332 6316
rect 371384 6304 371390 6316
rect 441522 6304 441528 6316
rect 371384 6276 441528 6304
rect 371384 6264 371390 6276
rect 441522 6264 441528 6276
rect 441580 6264 441586 6316
rect 234706 6196 234712 6248
rect 234764 6236 234770 6248
rect 305638 6236 305644 6248
rect 234764 6208 305644 6236
rect 234764 6196 234770 6208
rect 305638 6196 305644 6208
rect 305696 6196 305702 6248
rect 345014 6196 345020 6248
rect 345072 6236 345078 6248
rect 359918 6236 359924 6248
rect 345072 6208 359924 6236
rect 345072 6196 345078 6208
rect 359918 6196 359924 6208
rect 359976 6196 359982 6248
rect 371418 6196 371424 6248
rect 371476 6236 371482 6248
rect 445018 6236 445024 6248
rect 371476 6208 445024 6236
rect 371476 6196 371482 6208
rect 445018 6196 445024 6208
rect 445076 6196 445082 6248
rect 12342 6128 12348 6180
rect 12400 6168 12406 6180
rect 237742 6168 237748 6180
rect 12400 6140 237748 6168
rect 12400 6128 12406 6140
rect 237742 6128 237748 6140
rect 237800 6128 237806 6180
rect 242894 6128 242900 6180
rect 242952 6168 242958 6180
rect 302878 6168 302884 6180
rect 242952 6140 302884 6168
rect 242952 6128 242958 6140
rect 302878 6128 302884 6140
rect 302936 6128 302942 6180
rect 346486 6128 346492 6180
rect 346544 6168 346550 6180
rect 364610 6168 364616 6180
rect 346544 6140 364616 6168
rect 346544 6128 346550 6140
rect 364610 6128 364616 6140
rect 364668 6128 364674 6180
rect 412634 6128 412640 6180
rect 412692 6168 412698 6180
rect 576302 6168 576308 6180
rect 412692 6140 576308 6168
rect 412692 6128 412698 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 366358 5516 366364 5568
rect 366416 5556 366422 5568
rect 368198 5556 368204 5568
rect 366416 5528 368204 5556
rect 366416 5516 366422 5528
rect 368198 5516 368204 5528
rect 368256 5516 368262 5568
rect 303154 5176 303160 5228
rect 303212 5216 303218 5228
rect 328546 5216 328552 5228
rect 303212 5188 328552 5216
rect 303212 5176 303218 5188
rect 328546 5176 328552 5188
rect 328604 5176 328610 5228
rect 299658 5108 299664 5160
rect 299716 5148 299722 5160
rect 327350 5148 327356 5160
rect 299716 5120 327356 5148
rect 299716 5108 299722 5120
rect 327350 5108 327356 5120
rect 327408 5108 327414 5160
rect 296070 5040 296076 5092
rect 296128 5080 296134 5092
rect 325786 5080 325792 5092
rect 296128 5052 325792 5080
rect 296128 5040 296134 5052
rect 325786 5040 325792 5052
rect 325844 5040 325850 5092
rect 288986 4972 288992 5024
rect 289044 5012 289050 5024
rect 323026 5012 323032 5024
rect 289044 4984 323032 5012
rect 289044 4972 289050 4984
rect 323026 4972 323032 4984
rect 323084 4972 323090 5024
rect 285398 4904 285404 4956
rect 285456 4944 285462 4956
rect 323118 4944 323124 4956
rect 285456 4916 323124 4944
rect 285456 4904 285462 4916
rect 323118 4904 323124 4916
rect 323176 4904 323182 4956
rect 278314 4836 278320 4888
rect 278372 4876 278378 4888
rect 320358 4876 320364 4888
rect 278372 4848 320364 4876
rect 278372 4836 278378 4848
rect 320358 4836 320364 4848
rect 320416 4836 320422 4888
rect 351178 4836 351184 4888
rect 351236 4876 351242 4888
rect 356330 4876 356336 4888
rect 351236 4848 356336 4876
rect 351236 4836 351242 4848
rect 356330 4836 356336 4848
rect 356388 4836 356394 4888
rect 218146 4768 218152 4820
rect 218204 4808 218210 4820
rect 233878 4808 233884 4820
rect 218204 4780 233884 4808
rect 218204 4768 218210 4780
rect 233878 4768 233884 4780
rect 233936 4768 233942 4820
rect 246390 4768 246396 4820
rect 246448 4808 246454 4820
rect 289078 4808 289084 4820
rect 246448 4780 289084 4808
rect 246448 4768 246454 4780
rect 289078 4768 289084 4780
rect 289136 4768 289142 4820
rect 292574 4768 292580 4820
rect 292632 4808 292638 4820
rect 324498 4808 324504 4820
rect 292632 4780 324504 4808
rect 292632 4768 292638 4780
rect 324498 4768 324504 4780
rect 324556 4768 324562 4820
rect 354674 4768 354680 4820
rect 354732 4808 354738 4820
rect 391842 4808 391848 4820
rect 354732 4780 391848 4808
rect 354732 4768 354738 4780
rect 391842 4768 391848 4780
rect 391900 4768 391906 4820
rect 401594 4768 401600 4820
rect 401652 4808 401658 4820
rect 540790 4808 540796 4820
rect 401652 4780 540796 4808
rect 401652 4768 401658 4780
rect 540790 4768 540796 4780
rect 540848 4768 540854 4820
rect 382918 4496 382924 4548
rect 382976 4536 382982 4548
rect 384758 4536 384764 4548
rect 382976 4508 384764 4536
rect 382976 4496 382982 4508
rect 384758 4496 384764 4508
rect 384816 4496 384822 4548
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 176654 4156 176660 4208
rect 176712 4196 176718 4208
rect 177850 4196 177856 4208
rect 176712 4168 177856 4196
rect 176712 4156 176718 4168
rect 177850 4156 177856 4168
rect 177908 4156 177914 4208
rect 345658 4156 345664 4208
rect 345716 4196 345722 4208
rect 352834 4196 352840 4208
rect 345716 4168 352840 4196
rect 345716 4156 345722 4168
rect 352834 4156 352840 4168
rect 352892 4156 352898 4208
rect 103330 4088 103336 4140
rect 103388 4128 103394 4140
rect 266630 4128 266636 4140
rect 103388 4100 266636 4128
rect 103388 4088 103394 4100
rect 266630 4088 266636 4100
rect 266688 4088 266694 4140
rect 305546 4088 305552 4140
rect 305604 4128 305610 4140
rect 328454 4128 328460 4140
rect 305604 4100 328460 4128
rect 305604 4088 305610 4100
rect 328454 4088 328460 4100
rect 328512 4088 328518 4140
rect 333882 4088 333888 4140
rect 333940 4128 333946 4140
rect 336826 4128 336832 4140
rect 333940 4100 336832 4128
rect 333940 4088 333946 4100
rect 336826 4088 336832 4100
rect 336884 4088 336890 4140
rect 367094 4088 367100 4140
rect 367152 4128 367158 4140
rect 429654 4128 429660 4140
rect 367152 4100 429660 4128
rect 367152 4088 367158 4100
rect 429654 4088 429660 4100
rect 429712 4088 429718 4140
rect 46658 4020 46664 4072
rect 46716 4060 46722 4072
rect 248690 4060 248696 4072
rect 46716 4032 248696 4060
rect 46716 4020 46722 4032
rect 248690 4020 248696 4032
rect 248748 4020 248754 4072
rect 301958 4020 301964 4072
rect 302016 4060 302022 4072
rect 327258 4060 327264 4072
rect 302016 4032 327264 4060
rect 302016 4020 302022 4032
rect 327258 4020 327264 4032
rect 327316 4020 327322 4072
rect 332686 4020 332692 4072
rect 332744 4060 332750 4072
rect 337102 4060 337108 4072
rect 332744 4032 337108 4060
rect 332744 4020 332750 4032
rect 337102 4020 337108 4032
rect 337160 4020 337166 4072
rect 340874 4020 340880 4072
rect 340932 4060 340938 4072
rect 346946 4060 346952 4072
rect 340932 4032 346952 4060
rect 340932 4020 340938 4032
rect 346946 4020 346952 4032
rect 347004 4020 347010 4072
rect 368474 4020 368480 4072
rect 368532 4060 368538 4072
rect 433242 4060 433248 4072
rect 368532 4032 433248 4060
rect 368532 4020 368538 4032
rect 433242 4020 433248 4032
rect 433300 4020 433306 4072
rect 43070 3952 43076 4004
rect 43128 3992 43134 4004
rect 247034 3992 247040 4004
rect 43128 3964 247040 3992
rect 43128 3952 43134 3964
rect 247034 3952 247040 3964
rect 247092 3952 247098 4004
rect 298462 3952 298468 4004
rect 298520 3992 298526 4004
rect 327166 3992 327172 4004
rect 298520 3964 327172 3992
rect 298520 3952 298526 3964
rect 327166 3952 327172 3964
rect 327224 3952 327230 4004
rect 330386 3952 330392 4004
rect 330444 3992 330450 4004
rect 336918 3992 336924 4004
rect 330444 3964 336924 3992
rect 330444 3952 330450 3964
rect 336918 3952 336924 3964
rect 336976 3952 336982 4004
rect 368566 3952 368572 4004
rect 368624 3992 368630 4004
rect 436738 3992 436744 4004
rect 368624 3964 436744 3992
rect 368624 3952 368630 3964
rect 436738 3952 436744 3964
rect 436796 3952 436802 4004
rect 39574 3884 39580 3936
rect 39632 3924 39638 3936
rect 247126 3924 247132 3936
rect 39632 3896 247132 3924
rect 39632 3884 39638 3896
rect 247126 3884 247132 3896
rect 247184 3884 247190 3936
rect 294874 3884 294880 3936
rect 294932 3924 294938 3936
rect 325878 3924 325884 3936
rect 294932 3896 325884 3924
rect 294932 3884 294938 3896
rect 325878 3884 325884 3896
rect 325936 3884 325942 3936
rect 369854 3884 369860 3936
rect 369912 3924 369918 3936
rect 440326 3924 440332 3936
rect 369912 3896 440332 3924
rect 369912 3884 369918 3896
rect 440326 3884 440332 3896
rect 440384 3884 440390 3936
rect 35986 3816 35992 3868
rect 36044 3856 36050 3868
rect 245930 3856 245936 3868
rect 36044 3828 245936 3856
rect 36044 3816 36050 3828
rect 245930 3816 245936 3828
rect 245988 3816 245994 3868
rect 291378 3816 291384 3868
rect 291436 3856 291442 3868
rect 324406 3856 324412 3868
rect 291436 3828 324412 3856
rect 291436 3816 291442 3828
rect 324406 3816 324412 3828
rect 324464 3816 324470 3868
rect 329006 3816 329012 3868
rect 329064 3856 329070 3868
rect 334158 3856 334164 3868
rect 329064 3828 334164 3856
rect 329064 3816 329070 3828
rect 334158 3816 334164 3828
rect 334216 3816 334222 3868
rect 342622 3816 342628 3868
rect 342680 3856 342686 3868
rect 349246 3856 349252 3868
rect 342680 3828 349252 3856
rect 342680 3816 342686 3828
rect 349246 3816 349252 3828
rect 349304 3816 349310 3868
rect 371234 3816 371240 3868
rect 371292 3856 371298 3868
rect 443822 3856 443828 3868
rect 371292 3828 443828 3856
rect 371292 3816 371298 3828
rect 443822 3816 443828 3828
rect 443880 3816 443886 3868
rect 32398 3748 32404 3800
rect 32456 3788 32462 3800
rect 244274 3788 244280 3800
rect 32456 3760 244280 3788
rect 32456 3748 32462 3760
rect 244274 3748 244280 3760
rect 244332 3748 244338 3800
rect 287790 3748 287796 3800
rect 287848 3788 287854 3800
rect 322934 3788 322940 3800
rect 287848 3760 322940 3788
rect 287848 3748 287854 3760
rect 322934 3748 322940 3760
rect 322992 3748 322998 3800
rect 326798 3748 326804 3800
rect 326856 3788 326862 3800
rect 335446 3788 335452 3800
rect 326856 3760 335452 3788
rect 326856 3748 326862 3760
rect 335446 3748 335452 3760
rect 335504 3748 335510 3800
rect 342346 3748 342352 3800
rect 342404 3788 342410 3800
rect 348050 3788 348056 3800
rect 342404 3760 348056 3788
rect 342404 3748 342410 3760
rect 348050 3748 348056 3760
rect 348108 3748 348114 3800
rect 374178 3748 374184 3800
rect 374236 3788 374242 3800
rect 450906 3788 450912 3800
rect 374236 3760 450912 3788
rect 374236 3748 374242 3760
rect 450906 3748 450912 3760
rect 450964 3748 450970 3800
rect 576118 3748 576124 3800
rect 576176 3788 576182 3800
rect 578602 3788 578608 3800
rect 576176 3760 578608 3788
rect 576176 3748 576182 3760
rect 578602 3748 578608 3760
rect 578660 3748 578666 3800
rect 28902 3680 28908 3732
rect 28960 3720 28966 3732
rect 243170 3720 243176 3732
rect 28960 3692 243176 3720
rect 28960 3680 28966 3692
rect 243170 3680 243176 3692
rect 243228 3680 243234 3732
rect 284294 3680 284300 3732
rect 284352 3720 284358 3732
rect 321646 3720 321652 3732
rect 284352 3692 321652 3720
rect 284352 3680 284358 3692
rect 321646 3680 321652 3692
rect 321704 3680 321710 3732
rect 323302 3680 323308 3732
rect 323360 3720 323366 3732
rect 334066 3720 334072 3732
rect 323360 3692 334072 3720
rect 323360 3680 323366 3692
rect 334066 3680 334072 3692
rect 334124 3680 334130 3732
rect 342530 3680 342536 3732
rect 342588 3720 342594 3732
rect 350442 3720 350448 3732
rect 342588 3692 350448 3720
rect 342588 3680 342594 3692
rect 350442 3680 350448 3692
rect 350500 3680 350506 3732
rect 375374 3680 375380 3732
rect 375432 3720 375438 3732
rect 458082 3720 458088 3732
rect 375432 3692 458088 3720
rect 375432 3680 375438 3692
rect 458082 3680 458088 3692
rect 458140 3680 458146 3732
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 241606 3652 241612 3664
rect 25372 3624 241612 3652
rect 25372 3612 25378 3624
rect 241606 3612 241612 3624
rect 241664 3612 241670 3664
rect 280706 3612 280712 3664
rect 280764 3652 280770 3664
rect 321830 3652 321836 3664
rect 280764 3624 321836 3652
rect 280764 3612 280770 3624
rect 321830 3612 321836 3624
rect 321888 3612 321894 3664
rect 325602 3612 325608 3664
rect 325660 3652 325666 3664
rect 335538 3652 335544 3664
rect 325660 3624 335544 3652
rect 325660 3612 325666 3624
rect 335538 3612 335544 3624
rect 335596 3612 335602 3664
rect 346394 3612 346400 3664
rect 346452 3652 346458 3664
rect 362310 3652 362316 3664
rect 346452 3624 362316 3652
rect 346452 3612 346458 3624
rect 362310 3612 362316 3624
rect 362368 3612 362374 3664
rect 378134 3612 378140 3664
rect 378192 3652 378198 3664
rect 465166 3652 465172 3664
rect 378192 3624 465172 3652
rect 378192 3612 378198 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 241514 3584 241520 3596
rect 24268 3556 241520 3584
rect 24268 3544 24274 3556
rect 241514 3544 241520 3556
rect 241572 3544 241578 3596
rect 268010 3544 268016 3596
rect 268068 3584 268074 3596
rect 268470 3584 268476 3596
rect 268068 3556 268476 3584
rect 268068 3544 268074 3556
rect 268470 3544 268476 3556
rect 268528 3544 268534 3596
rect 271874 3544 271880 3596
rect 271932 3584 271938 3596
rect 272058 3584 272064 3596
rect 271932 3556 272064 3584
rect 271932 3544 271938 3556
rect 272058 3544 272064 3556
rect 272116 3544 272122 3596
rect 273622 3544 273628 3596
rect 273680 3584 273686 3596
rect 318794 3584 318800 3596
rect 273680 3556 318800 3584
rect 273680 3544 273686 3556
rect 318794 3544 318800 3556
rect 318852 3544 318858 3596
rect 322106 3544 322112 3596
rect 322164 3584 322170 3596
rect 329006 3584 329012 3596
rect 322164 3556 329012 3584
rect 322164 3544 322170 3556
rect 329006 3544 329012 3556
rect 329064 3544 329070 3596
rect 332594 3584 332600 3596
rect 329116 3556 332600 3584
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6178 3516 6184 3528
rect 5316 3488 6184 3516
rect 5316 3476 5322 3488
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 10318 3516 10324 3528
rect 6288 3488 10324 3516
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 6288 3448 6316 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 15838 3516 15844 3528
rect 11204 3488 15844 3516
rect 11204 3476 11210 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 24118 3516 24124 3528
rect 18288 3488 24124 3516
rect 18288 3476 18294 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 240410 3516 240416 3528
rect 24320 3488 240416 3516
rect 4120 3420 6316 3448
rect 4120 3408 4126 3420
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 11698 3380 11704 3392
rect 1728 3352 11704 3380
rect 1728 3340 1734 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 24320 3380 24348 3488
rect 240410 3476 240416 3488
rect 240468 3476 240474 3528
rect 270034 3476 270040 3528
rect 270092 3516 270098 3528
rect 317690 3516 317696 3528
rect 270092 3488 317696 3516
rect 270092 3476 270098 3488
rect 317690 3476 317696 3488
rect 317748 3476 317754 3528
rect 319714 3476 319720 3528
rect 319772 3516 319778 3528
rect 329116 3516 329144 3556
rect 332594 3544 332600 3556
rect 332652 3544 332658 3596
rect 342438 3544 342444 3596
rect 342496 3584 342502 3596
rect 351638 3584 351644 3596
rect 342496 3556 351644 3584
rect 342496 3544 342502 3556
rect 351638 3544 351644 3556
rect 351696 3544 351702 3596
rect 360194 3544 360200 3596
rect 360252 3584 360258 3596
rect 408402 3584 408408 3596
rect 360252 3556 408408 3584
rect 360252 3544 360258 3556
rect 408402 3544 408408 3556
rect 408460 3544 408466 3596
rect 414106 3544 414112 3596
rect 414164 3584 414170 3596
rect 580994 3584 581000 3596
rect 414164 3556 581000 3584
rect 414164 3544 414170 3556
rect 580994 3544 581000 3556
rect 581052 3544 581058 3596
rect 319772 3488 329144 3516
rect 319772 3476 319778 3488
rect 331582 3476 331588 3528
rect 331640 3516 331646 3528
rect 333238 3516 333244 3528
rect 331640 3488 333244 3516
rect 331640 3476 331646 3488
rect 333238 3476 333244 3488
rect 333296 3476 333302 3528
rect 337470 3476 337476 3528
rect 337528 3516 337534 3528
rect 338390 3516 338396 3528
rect 337528 3488 338396 3516
rect 337528 3476 337534 3488
rect 338390 3476 338396 3488
rect 338448 3476 338454 3528
rect 338666 3476 338672 3528
rect 338724 3516 338730 3528
rect 339586 3516 339592 3528
rect 338724 3488 339592 3516
rect 338724 3476 338730 3488
rect 339586 3476 339592 3488
rect 339644 3476 339650 3528
rect 339678 3476 339684 3528
rect 339736 3516 339742 3528
rect 340966 3516 340972 3528
rect 339736 3488 340972 3516
rect 339736 3476 339742 3488
rect 340966 3476 340972 3488
rect 341024 3476 341030 3528
rect 343634 3476 343640 3528
rect 343692 3516 343698 3528
rect 354030 3516 354036 3528
rect 343692 3488 354036 3516
rect 343692 3476 343698 3488
rect 354030 3476 354036 3488
rect 354088 3476 354094 3528
rect 357434 3476 357440 3528
rect 357492 3516 357498 3528
rect 358722 3516 358728 3528
rect 357492 3488 358728 3516
rect 357492 3476 357498 3488
rect 358722 3476 358728 3488
rect 358780 3476 358786 3528
rect 373994 3476 374000 3528
rect 374052 3516 374058 3528
rect 375282 3516 375288 3528
rect 374052 3488 375288 3516
rect 374052 3476 374058 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 379514 3476 379520 3528
rect 379572 3516 379578 3528
rect 472250 3516 472256 3528
rect 379572 3488 472256 3516
rect 379572 3476 379578 3488
rect 472250 3476 472256 3488
rect 472308 3476 472314 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 240226 3448 240232 3460
rect 20680 3352 24348 3380
rect 26206 3420 240232 3448
rect 20680 3340 20686 3352
rect 13538 3272 13544 3324
rect 13596 3312 13602 3324
rect 18598 3312 18604 3324
rect 13596 3284 18604 3312
rect 13596 3272 13602 3284
rect 18598 3272 18604 3284
rect 18656 3272 18662 3324
rect 19426 3272 19432 3324
rect 19484 3312 19490 3324
rect 26206 3312 26234 3420
rect 240226 3408 240232 3420
rect 240284 3408 240290 3460
rect 266538 3408 266544 3460
rect 266596 3448 266602 3460
rect 316034 3448 316040 3460
rect 266596 3420 316040 3448
rect 266596 3408 266602 3420
rect 316034 3408 316040 3420
rect 316092 3408 316098 3460
rect 318518 3408 318524 3460
rect 318576 3448 318582 3460
rect 332778 3448 332784 3460
rect 318576 3420 332784 3448
rect 318576 3408 318582 3420
rect 332778 3408 332784 3420
rect 332836 3408 332842 3460
rect 343726 3408 343732 3460
rect 343784 3448 343790 3460
rect 355226 3448 355232 3460
rect 343784 3420 355232 3448
rect 343784 3408 343790 3420
rect 355226 3408 355232 3420
rect 355284 3408 355290 3460
rect 361574 3408 361580 3460
rect 361632 3448 361638 3460
rect 411898 3448 411904 3460
rect 361632 3420 411904 3448
rect 361632 3408 361638 3420
rect 411898 3408 411904 3420
rect 411956 3408 411962 3460
rect 415394 3408 415400 3460
rect 415452 3448 415458 3460
rect 416682 3448 416688 3460
rect 415452 3420 416688 3448
rect 415452 3408 415458 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 416774 3408 416780 3460
rect 416832 3448 416838 3460
rect 582190 3448 582196 3460
rect 416832 3420 582196 3448
rect 416832 3408 416838 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 77294 3340 77300 3392
rect 77352 3380 77358 3392
rect 78214 3380 78220 3392
rect 77352 3352 78220 3380
rect 77352 3340 77358 3352
rect 78214 3340 78220 3352
rect 78272 3340 78278 3392
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 106918 3340 106924 3392
rect 106976 3380 106982 3392
rect 268194 3380 268200 3392
rect 106976 3352 268200 3380
rect 106976 3340 106982 3352
rect 268194 3340 268200 3352
rect 268252 3340 268258 3392
rect 309042 3340 309048 3392
rect 309100 3380 309106 3392
rect 329834 3380 329840 3392
rect 309100 3352 329840 3380
rect 309100 3340 309106 3352
rect 329834 3340 329840 3352
rect 329892 3340 329898 3392
rect 341058 3340 341064 3392
rect 341116 3380 341122 3392
rect 344554 3380 344560 3392
rect 341116 3352 344560 3380
rect 341116 3340 341122 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 426158 3380 426164 3392
rect 365772 3352 426164 3380
rect 365772 3340 365778 3352
rect 426158 3340 426164 3352
rect 426216 3340 426222 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 19484 3284 26234 3312
rect 19484 3272 19490 3284
rect 118694 3272 118700 3324
rect 118752 3312 118758 3324
rect 119890 3312 119896 3324
rect 118752 3284 119896 3312
rect 118752 3272 118758 3284
rect 119890 3272 119896 3284
rect 119948 3272 119954 3324
rect 269114 3312 269120 3324
rect 120000 3284 269120 3312
rect 9950 3204 9956 3256
rect 10008 3244 10014 3256
rect 13170 3244 13176 3256
rect 10008 3216 13176 3244
rect 10008 3204 10014 3216
rect 13170 3204 13176 3216
rect 13228 3204 13234 3256
rect 114002 3204 114008 3256
rect 114060 3244 114066 3256
rect 120000 3244 120028 3284
rect 269114 3272 269120 3284
rect 269172 3272 269178 3324
rect 312630 3272 312636 3324
rect 312688 3312 312694 3324
rect 331398 3312 331404 3324
rect 312688 3284 331404 3312
rect 312688 3272 312694 3284
rect 331398 3272 331404 3284
rect 331456 3272 331462 3324
rect 364426 3272 364432 3324
rect 364484 3312 364490 3324
rect 422570 3312 422576 3324
rect 364484 3284 422576 3312
rect 364484 3272 364490 3284
rect 422570 3272 422576 3284
rect 422628 3272 422634 3324
rect 114060 3216 120028 3244
rect 114060 3204 114066 3216
rect 121086 3204 121092 3256
rect 121144 3244 121150 3256
rect 271874 3244 271880 3256
rect 121144 3216 271880 3244
rect 121144 3204 121150 3216
rect 271874 3204 271880 3216
rect 271932 3204 271938 3256
rect 315022 3204 315028 3256
rect 315080 3244 315086 3256
rect 331214 3244 331220 3256
rect 315080 3216 331220 3244
rect 315080 3204 315086 3216
rect 331214 3204 331220 3216
rect 331272 3204 331278 3256
rect 364334 3204 364340 3256
rect 364392 3244 364398 3256
rect 418982 3244 418988 3256
rect 364392 3216 418988 3244
rect 364392 3204 364398 3216
rect 418982 3204 418988 3216
rect 419040 3204 419046 3256
rect 23014 3136 23020 3188
rect 23072 3176 23078 3188
rect 25498 3176 25504 3188
rect 23072 3148 25504 3176
rect 23072 3136 23078 3148
rect 25498 3136 25504 3148
rect 25556 3136 25562 3188
rect 218054 3136 218060 3188
rect 218112 3176 218118 3188
rect 219250 3176 219256 3188
rect 218112 3148 219256 3176
rect 218112 3136 218118 3148
rect 219250 3136 219256 3148
rect 219308 3136 219314 3188
rect 234614 3136 234620 3188
rect 234672 3176 234678 3188
rect 235810 3176 235816 3188
rect 234672 3148 235816 3176
rect 234672 3136 234678 3148
rect 235810 3136 235816 3148
rect 235868 3136 235874 3188
rect 316218 3136 316224 3188
rect 316276 3176 316282 3188
rect 331306 3176 331312 3188
rect 316276 3148 331312 3176
rect 316276 3136 316282 3148
rect 331306 3136 331312 3148
rect 331364 3136 331370 3188
rect 336274 3136 336280 3188
rect 336332 3176 336338 3188
rect 338206 3176 338212 3188
rect 336332 3148 338212 3176
rect 336332 3136 336338 3148
rect 338206 3136 338212 3148
rect 338264 3136 338270 3188
rect 398926 3136 398932 3188
rect 398984 3176 398990 3188
rect 400122 3176 400128 3188
rect 398984 3148 400128 3176
rect 398984 3136 398990 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 414014 3136 414020 3188
rect 414072 3176 414078 3188
rect 416774 3176 416780 3188
rect 414072 3148 416780 3176
rect 414072 3136 414078 3148
rect 416774 3136 416780 3148
rect 416832 3136 416838 3188
rect 566 3068 572 3120
rect 624 3108 630 3120
rect 4798 3108 4804 3120
rect 624 3080 4804 3108
rect 624 3068 630 3080
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 329190 3000 329196 3052
rect 329248 3040 329254 3052
rect 335630 3040 335636 3052
rect 329248 3012 335636 3040
rect 329248 3000 329254 3012
rect 335630 3000 335636 3012
rect 335688 3000 335694 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 341150 2864 341156 2916
rect 341208 2904 341214 2916
rect 345750 2904 345756 2916
rect 341208 2876 345756 2904
rect 341208 2864 341214 2876
rect 345750 2864 345756 2876
rect 345808 2864 345814 2916
rect 299474 2048 299480 2100
rect 299532 2088 299538 2100
rect 300762 2088 300768 2100
rect 299532 2060 300768 2088
rect 299532 2048 299538 2060
rect 300762 2048 300768 2060
rect 300820 2048 300826 2100
rect 423674 960 423680 1012
rect 423732 1000 423738 1012
rect 424962 1000 424968 1012
rect 423732 972 424968 1000
rect 423732 960 423738 972
rect 424962 960 424968 972
rect 425020 960 425026 1012
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 283840 700748 283892 700800
rect 328460 700748 328512 700800
rect 318800 700680 318852 700732
rect 413652 700680 413704 700732
rect 218980 700612 219032 700664
rect 332600 700612 332652 700664
rect 154120 700544 154172 700596
rect 338120 700544 338172 700596
rect 89168 700476 89220 700528
rect 342260 700476 342312 700528
rect 72976 700408 73028 700460
rect 340880 700408 340932 700460
rect 24308 700340 24360 700392
rect 347872 700340 347924 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 460204 700272 460256 700324
rect 559656 700272 559708 700324
rect 235172 698912 235224 698964
rect 329840 698912 329892 698964
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 303620 696940 303672 696992
rect 580172 696940 580224 696992
rect 305000 683136 305052 683188
rect 580172 683136 580224 683188
rect 300860 670760 300912 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 351920 670692 351972 670744
rect 306380 660288 306432 660340
rect 460204 660288 460256 660340
rect 3516 656888 3568 656940
rect 350540 656888 350592 656940
rect 298100 643084 298152 643136
rect 580172 643084 580224 643136
rect 299572 630640 299624 630692
rect 580172 630640 580224 630692
rect 3332 618264 3384 618316
rect 356060 618264 356112 618316
rect 296720 616836 296772 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 354680 605820 354732 605872
rect 293960 590656 294012 590708
rect 579804 590656 579856 590708
rect 295340 576852 295392 576904
rect 580172 576852 580224 576904
rect 3056 565836 3108 565888
rect 361580 565836 361632 565888
rect 292580 563048 292632 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 360200 553392 360252 553444
rect 288440 536800 288492 536852
rect 580172 536800 580224 536852
rect 320180 527824 320232 527876
rect 364340 527824 364392 527876
rect 289820 524424 289872 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 365720 514768 365772 514820
rect 287060 510620 287112 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 364340 500964 364392 501016
rect 284300 484372 284352 484424
rect 580172 484372 580224 484424
rect 285864 470568 285916 470620
rect 579988 470568 580040 470620
rect 104900 468460 104952 468512
rect 339592 468460 339644 468512
rect 169760 467100 169812 467152
rect 334808 467100 334860 467152
rect 299480 465672 299532 465724
rect 325700 465672 325752 465724
rect 316040 464312 316092 464364
rect 429200 464312 429252 464364
rect 226984 462476 227036 462528
rect 375932 462476 375984 462528
rect 225604 462408 225656 462460
rect 380900 462408 380952 462460
rect 3516 462340 3568 462392
rect 371240 462340 371292 462392
rect 311808 461592 311860 461644
rect 494060 461592 494112 461644
rect 233976 461320 234028 461372
rect 369860 461320 369912 461372
rect 280068 461252 280120 461304
rect 417516 461252 417568 461304
rect 278688 461184 278740 461236
rect 422944 461184 422996 461236
rect 273996 461116 274048 461168
rect 420184 461116 420236 461168
rect 228364 461048 228416 461100
rect 379152 461048 379204 461100
rect 229744 460980 229796 461032
rect 396540 460980 396592 461032
rect 4896 460912 4948 460964
rect 391940 460912 391992 460964
rect 318156 460844 318208 460896
rect 397460 460844 397512 460896
rect 201500 460776 201552 460828
rect 331772 460776 331824 460828
rect 313096 460708 313148 460760
rect 462320 460708 462372 460760
rect 315028 460640 315080 460692
rect 477500 460640 477552 460692
rect 136640 460572 136692 460624
rect 336740 460572 336792 460624
rect 308680 460504 308732 460556
rect 527180 460504 527232 460556
rect 310244 460436 310296 460488
rect 542360 460436 542412 460488
rect 3608 460368 3660 460420
rect 353852 460368 353904 460420
rect 3700 460300 3752 460352
rect 358820 460300 358872 460352
rect 3792 460232 3844 460284
rect 363328 460232 363380 460284
rect 3884 460164 3936 460216
rect 368112 460164 368164 460216
rect 266360 460096 266412 460148
rect 327080 460096 327132 460148
rect 324136 460028 324188 460080
rect 347780 460028 347832 460080
rect 322848 459960 322900 460012
rect 331220 459960 331272 460012
rect 355968 459552 356020 459604
rect 374368 459552 374420 459604
rect 233884 458804 233936 458856
rect 377588 458804 377640 458856
rect 275560 458736 275612 458788
rect 424324 458736 424376 458788
rect 277124 458668 277176 458720
rect 425704 458668 425756 458720
rect 232504 458600 232556 458652
rect 382280 458600 382332 458652
rect 231124 458532 231176 458584
rect 387064 458532 387116 458584
rect 255044 458464 255096 458516
rect 421564 458464 421616 458516
rect 245568 458396 245620 458448
rect 418804 458396 418856 458448
rect 240784 458328 240836 458380
rect 417424 458328 417476 458380
rect 235908 458260 235960 458312
rect 580264 458260 580316 458312
rect 3516 458192 3568 458244
rect 373126 458192 373178 458244
rect 3424 457444 3476 457496
rect 281632 457580 281684 457632
rect 283380 457444 283432 457496
rect 355968 457444 356020 457496
rect 427084 456832 427136 456884
rect 580172 456764 580224 456816
rect 3332 449828 3384 449880
rect 233976 449828 234028 449880
rect 417516 431876 417568 431928
rect 580172 431876 580224 431928
rect 427084 419432 427136 419484
rect 580172 419432 580224 419484
rect 2964 411204 3016 411256
rect 226984 411204 227036 411256
rect 422944 405628 422996 405680
rect 579620 405628 579672 405680
rect 424324 379448 424376 379500
rect 580172 379448 580224 379500
rect 3240 372512 3292 372564
rect 233884 372512 233936 372564
rect 425704 365644 425756 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 225604 358708 225656 358760
rect 420184 353200 420236 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 228364 346332 228416 346384
rect 294420 336744 294472 336796
rect 233976 336676 234028 336728
rect 237012 336676 237064 336728
rect 239404 336676 239456 336728
rect 240140 336676 240192 336728
rect 260840 336676 260892 336728
rect 261116 336676 261168 336728
rect 271144 336676 271196 336728
rect 272432 336676 272484 336728
rect 293224 336676 293276 336728
rect 296812 336676 296864 336728
rect 297272 336676 297324 336728
rect 300768 336676 300820 336728
rect 304080 336676 304132 336728
rect 309324 336676 309376 336728
rect 309508 336676 309560 336728
rect 335452 336676 335504 336728
rect 335636 336676 335688 336728
rect 346400 336676 346452 336728
rect 346676 336676 346728 336728
rect 367100 336676 367152 336728
rect 367468 336676 367520 336728
rect 376760 336676 376812 336728
rect 377036 336676 377088 336728
rect 386420 336676 386472 336728
rect 386788 336676 386840 336728
rect 397552 336676 397604 336728
rect 397828 336676 397880 336728
rect 401600 336676 401652 336728
rect 401876 336676 401928 336728
rect 367192 336608 367244 336660
rect 367744 336608 367796 336660
rect 253204 336540 253256 336592
rect 253940 336540 253992 336592
rect 289176 336540 289228 336592
rect 290004 336540 290056 336592
rect 298744 336540 298796 336592
rect 302424 336540 302476 336592
rect 340788 336540 340840 336592
rect 341340 336540 341392 336592
rect 399760 336540 399812 336592
rect 400864 336540 400916 336592
rect 269764 336472 269816 336524
rect 271880 336472 271932 336524
rect 294604 336472 294656 336524
rect 298560 336472 298612 336524
rect 303068 336472 303120 336524
rect 305368 336472 305420 336524
rect 350080 336472 350132 336524
rect 358084 336472 358136 336524
rect 362868 336472 362920 336524
rect 373356 336472 373408 336524
rect 233884 336404 233936 336456
rect 124220 336336 124272 336388
rect 273260 336336 273312 336388
rect 297456 336404 297508 336456
rect 299848 336404 299900 336456
rect 302884 336404 302936 336456
rect 309692 336404 309744 336456
rect 353760 336404 353812 336456
rect 382924 336404 382976 336456
rect 302240 336336 302292 336388
rect 305828 336336 305880 336388
rect 313372 336336 313424 336388
rect 358176 336336 358228 336388
rect 387064 336336 387116 336388
rect 396448 336336 396500 336388
rect 422944 336336 422996 336388
rect 117320 336268 117372 336320
rect 271052 336268 271104 336320
rect 286416 336268 286468 336320
rect 287796 336268 287848 336320
rect 302976 336268 303028 336320
rect 314844 336268 314896 336320
rect 315304 336268 315356 336320
rect 324320 336268 324372 336320
rect 334348 336268 334400 336320
rect 338212 336268 338264 336320
rect 343824 336268 343876 336320
rect 345664 336268 345716 336320
rect 345756 336268 345808 336320
rect 357440 336268 357492 336320
rect 362776 336268 362828 336320
rect 370504 336268 370556 336320
rect 373080 336268 373132 336320
rect 447140 336268 447192 336320
rect 110420 336200 110472 336252
rect 268844 336200 268896 336252
rect 307024 336200 307076 336252
rect 322112 336200 322164 336252
rect 339500 336200 339552 336252
rect 339684 336200 339736 336252
rect 347320 336200 347372 336252
rect 362960 336200 363012 336252
rect 375288 336200 375340 336252
rect 454040 336200 454092 336252
rect 99380 336132 99432 336184
rect 265532 336132 265584 336184
rect 297364 336132 297416 336184
rect 311900 336132 311952 336184
rect 324320 336132 324372 336184
rect 334900 336132 334952 336184
rect 348608 336132 348660 336184
rect 359464 336132 359516 336184
rect 377496 336132 377548 336184
rect 460940 336132 460992 336184
rect 15844 336064 15896 336116
rect 238116 336064 238168 336116
rect 276664 336064 276716 336116
rect 285680 336064 285732 336116
rect 289084 336064 289136 336116
rect 310796 336064 310848 336116
rect 327080 336064 327132 336116
rect 336004 336064 336056 336116
rect 350816 336064 350868 336116
rect 374000 336064 374052 336116
rect 379888 336064 379940 336116
rect 467840 336064 467892 336116
rect 6184 335996 6236 336048
rect 236276 335996 236328 336048
rect 269304 335996 269356 336048
rect 284484 335996 284536 336048
rect 286232 335996 286284 336048
rect 291200 335996 291252 336048
rect 264244 335928 264296 335980
rect 267004 335928 267056 335980
rect 291844 335928 291896 335980
rect 315212 335996 315264 336048
rect 320180 335996 320232 336048
rect 333980 335996 334032 336048
rect 344928 335996 344980 336048
rect 351184 335996 351236 336048
rect 351920 335996 351972 336048
rect 377404 335996 377456 336048
rect 381820 335996 381872 336048
rect 474740 335996 474792 336048
rect 305644 335928 305696 335980
rect 307208 335928 307260 335980
rect 359464 335928 359516 335980
rect 366180 335928 366232 335980
rect 251824 335860 251876 335912
rect 253020 335860 253072 335912
rect 291936 335792 291988 335844
rect 293316 335792 293368 335844
rect 319444 335792 319496 335844
rect 321008 335792 321060 335844
rect 273904 335724 273956 335776
rect 277952 335724 278004 335776
rect 287704 335656 287756 335708
rect 290372 335656 290424 335708
rect 322204 335656 322256 335708
rect 326528 335656 326580 335708
rect 340972 335656 341024 335708
rect 342260 335656 342312 335708
rect 244924 335520 244976 335572
rect 246212 335520 246264 335572
rect 301504 335452 301556 335504
rect 308588 335452 308640 335504
rect 320824 335452 320876 335504
rect 327632 335452 327684 335504
rect 361764 335452 361816 335504
rect 364984 335452 365036 335504
rect 379980 335384 380032 335436
rect 381544 335384 381596 335436
rect 295984 335316 296036 335368
rect 296720 335316 296772 335368
rect 304264 335316 304316 335368
rect 307852 335316 307904 335368
rect 313924 335316 313976 335368
rect 317420 335316 317472 335368
rect 333244 335316 333296 335368
rect 337108 335316 337160 335368
rect 402336 335316 402388 335368
rect 403624 335316 403676 335368
rect 411812 335316 411864 335368
rect 413376 335316 413428 335368
rect 321652 335180 321704 335232
rect 321836 335180 321888 335232
rect 383568 334636 383620 334688
rect 480260 334636 480312 334688
rect 224960 334568 225012 334620
rect 300768 334568 300820 334620
rect 403164 334568 403216 334620
rect 543740 334568 543792 334620
rect 414020 334500 414072 334552
rect 414204 334500 414256 334552
rect 384488 333276 384540 333328
rect 483020 333276 483072 333328
rect 227720 333208 227772 333260
rect 303068 333208 303120 333260
rect 408500 333208 408552 333260
rect 561680 333208 561732 333260
rect 175280 331916 175332 331968
rect 288900 331916 288952 331968
rect 390008 331916 390060 331968
rect 500960 331916 501012 331968
rect 46940 331848 46992 331900
rect 249432 331848 249484 331900
rect 403808 331848 403860 331900
rect 546500 331848 546552 331900
rect 383844 331168 383896 331220
rect 384028 331168 384080 331220
rect 347964 330760 348016 330812
rect 238760 330624 238812 330676
rect 239588 330624 239640 330676
rect 168380 330556 168432 330608
rect 286692 330556 286744 330608
rect 347964 330556 348016 330608
rect 366272 330556 366324 330608
rect 423680 330556 423732 330608
rect 57980 330488 58032 330540
rect 234620 330420 234672 330472
rect 235540 330420 235592 330472
rect 238852 330488 238904 330540
rect 239220 330488 239272 330540
rect 240232 330488 240284 330540
rect 240692 330488 240744 330540
rect 241520 330488 241572 330540
rect 242164 330488 242216 330540
rect 243084 330488 243136 330540
rect 244004 330488 244056 330540
rect 254124 330488 254176 330540
rect 254952 330488 255004 330540
rect 255412 330488 255464 330540
rect 255688 330488 255740 330540
rect 256700 330488 256752 330540
rect 257160 330488 257212 330540
rect 258172 330488 258224 330540
rect 258632 330488 258684 330540
rect 259460 330488 259512 330540
rect 260380 330488 260432 330540
rect 260932 330488 260984 330540
rect 261852 330488 261904 330540
rect 262220 330488 262272 330540
rect 262956 330488 263008 330540
rect 265072 330488 265124 330540
rect 265900 330488 265952 330540
rect 266452 330488 266504 330540
rect 267372 330488 267424 330540
rect 267832 330488 267884 330540
rect 268292 330488 268344 330540
rect 269120 330488 269172 330540
rect 269948 330488 270000 330540
rect 270776 330488 270828 330540
rect 271328 330488 271380 330540
rect 271972 330488 272024 330540
rect 272800 330488 272852 330540
rect 285772 330488 285824 330540
rect 286324 330488 286376 330540
rect 291384 330488 291436 330540
rect 292212 330488 292264 330540
rect 302332 330488 302384 330540
rect 303160 330488 303212 330540
rect 305092 330488 305144 330540
rect 305736 330488 305788 330540
rect 306656 330488 306708 330540
rect 307484 330488 307536 330540
rect 309232 330488 309284 330540
rect 310060 330488 310112 330540
rect 310612 330488 310664 330540
rect 311164 330488 311216 330540
rect 313372 330488 313424 330540
rect 314108 330488 314160 330540
rect 314844 330488 314896 330540
rect 315580 330488 315632 330540
rect 316224 330488 316276 330540
rect 316684 330488 316736 330540
rect 318800 330488 318852 330540
rect 319260 330488 319312 330540
rect 331220 330488 331272 330540
rect 331956 330488 332008 330540
rect 332600 330488 332652 330540
rect 333428 330488 333480 330540
rect 334072 330488 334124 330540
rect 334532 330488 334584 330540
rect 336832 330488 336884 330540
rect 337844 330488 337896 330540
rect 342536 330488 342588 330540
rect 342996 330488 343048 330540
rect 345020 330488 345072 330540
rect 345848 330488 345900 330540
rect 347872 330488 347924 330540
rect 348792 330488 348844 330540
rect 360200 330488 360252 330540
rect 360844 330488 360896 330540
rect 364432 330488 364484 330540
rect 365260 330488 365312 330540
rect 367284 330488 367336 330540
rect 368112 330488 368164 330540
rect 368572 330488 368624 330540
rect 369584 330488 369636 330540
rect 390744 330488 390796 330540
rect 391204 330488 391256 330540
rect 392032 330488 392084 330540
rect 392584 330488 392636 330540
rect 393412 330488 393464 330540
rect 394424 330488 394476 330540
rect 396080 330488 396132 330540
rect 396632 330488 396684 330540
rect 397644 330488 397696 330540
rect 398472 330488 398524 330540
rect 255320 330420 255372 330472
rect 256424 330420 256476 330472
rect 256792 330420 256844 330472
rect 257528 330420 257580 330472
rect 258264 330420 258316 330472
rect 259000 330420 259052 330472
rect 262312 330420 262364 330472
rect 263324 330420 263376 330472
rect 316040 330420 316092 330472
rect 317052 330420 317104 330472
rect 331312 330420 331364 330472
rect 332324 330420 332376 330472
rect 342444 330420 342496 330472
rect 343272 330420 343324 330472
rect 390560 330420 390612 330472
rect 391480 330420 391532 330472
rect 391940 330420 391992 330472
rect 392952 330420 393004 330472
rect 396172 330420 396224 330472
rect 397000 330420 397052 330472
rect 397460 330420 397512 330472
rect 398104 330420 398156 330472
rect 252744 330352 252796 330404
rect 405280 330352 405332 330404
rect 550640 330488 550692 330540
rect 258080 330284 258132 330336
rect 258448 330284 258500 330336
rect 317512 330284 317564 330336
rect 318524 330284 318576 330336
rect 287152 330080 287204 330132
rect 288164 330080 288216 330132
rect 394700 329876 394752 329928
rect 395160 329876 395212 329928
rect 340972 329808 341024 329860
rect 341892 329808 341944 329860
rect 241612 329672 241664 329724
rect 242532 329672 242584 329724
rect 267924 329672 267976 329724
rect 268476 329672 268528 329724
rect 365812 329536 365864 329588
rect 366732 329536 366784 329588
rect 201500 329196 201552 329248
rect 296904 329196 296956 329248
rect 160100 329128 160152 329180
rect 269304 329128 269356 329180
rect 26240 329060 26292 329112
rect 242900 329060 242952 329112
rect 392124 329060 392176 329112
rect 507860 329060 507912 329112
rect 282920 328244 282972 328296
rect 283196 328244 283248 328296
rect 318984 328176 319036 328228
rect 319904 328176 319956 328228
rect 215300 327768 215352 327820
rect 301320 327768 301372 327820
rect 346492 327768 346544 327820
rect 347412 327768 347464 327820
rect 125600 327700 125652 327752
rect 273444 327700 273496 327752
rect 394056 327700 394108 327752
rect 514760 327700 514812 327752
rect 365720 327632 365772 327684
rect 366364 327632 366416 327684
rect 393320 327564 393372 327616
rect 393688 327564 393740 327616
rect 332692 327496 332744 327548
rect 333060 327496 333112 327548
rect 283012 326884 283064 326936
rect 283748 326884 283800 326936
rect 378324 326680 378376 326732
rect 280436 326476 280488 326528
rect 280620 326476 280672 326528
rect 354956 326476 355008 326528
rect 355140 326476 355192 326528
rect 375564 326476 375616 326528
rect 375748 326476 375800 326528
rect 378324 326476 378376 326528
rect 410064 326476 410116 326528
rect 410340 326476 410392 326528
rect 193220 326408 193272 326460
rect 293224 326408 293276 326460
rect 295524 326408 295576 326460
rect 323032 326408 323084 326460
rect 323952 326408 324004 326460
rect 328460 326408 328512 326460
rect 329104 326408 329156 326460
rect 354680 326408 354732 326460
rect 355692 326408 355744 326460
rect 356244 326408 356296 326460
rect 356428 326408 356480 326460
rect 371240 326408 371292 326460
rect 371792 326408 371844 326460
rect 372620 326408 372672 326460
rect 373632 326408 373684 326460
rect 374184 326408 374236 326460
rect 374736 326408 374788 326460
rect 375380 326408 375432 326460
rect 376208 326408 376260 326460
rect 376852 326408 376904 326460
rect 377680 326408 377732 326460
rect 378232 326408 378284 326460
rect 379152 326408 379204 326460
rect 379520 326408 379572 326460
rect 380532 326408 380584 326460
rect 381084 326408 381136 326460
rect 381268 326408 381320 326460
rect 382280 326408 382332 326460
rect 382740 326408 382792 326460
rect 383752 326408 383804 326460
rect 384580 326408 384632 326460
rect 385224 326408 385276 326460
rect 385684 326408 385736 326460
rect 386512 326408 386564 326460
rect 387156 326408 387208 326460
rect 387800 326408 387852 326460
rect 388628 326408 388680 326460
rect 398932 326408 398984 326460
rect 399116 326408 399168 326460
rect 401692 326408 401744 326460
rect 402520 326408 402572 326460
rect 403072 326408 403124 326460
rect 403900 326408 403952 326460
rect 404452 326408 404504 326460
rect 404636 326408 404688 326460
rect 405924 326408 405976 326460
rect 406476 326408 406528 326460
rect 407120 326408 407172 326460
rect 407580 326408 407632 326460
rect 409880 326408 409932 326460
rect 410524 326408 410576 326460
rect 411352 326408 411404 326460
rect 412364 326408 412416 326460
rect 4804 326340 4856 326392
rect 234804 326340 234856 326392
rect 244280 326340 244332 326392
rect 244740 326340 244792 326392
rect 245752 326340 245804 326392
rect 246580 326340 246632 326392
rect 247040 326340 247092 326392
rect 247960 326340 248012 326392
rect 249800 326340 249852 326392
rect 250168 326340 250220 326392
rect 251180 326340 251232 326392
rect 252008 326340 252060 326392
rect 273352 326340 273404 326392
rect 274272 326340 274324 326392
rect 274640 326340 274692 326392
rect 275008 326340 275060 326392
rect 276020 326340 276072 326392
rect 276480 326340 276532 326392
rect 277492 326340 277544 326392
rect 278320 326340 278372 326392
rect 278964 326340 279016 326392
rect 279424 326340 279476 326392
rect 280252 326340 280304 326392
rect 281264 326340 281316 326392
rect 281540 326340 281592 326392
rect 282000 326340 282052 326392
rect 294236 326340 294288 326392
rect 295156 326340 295208 326392
rect 249892 326272 249944 326324
rect 250904 326272 250956 326324
rect 278780 326272 278832 326324
rect 279792 326272 279844 326324
rect 296996 326340 297048 326392
rect 297640 326340 297692 326392
rect 299572 326340 299624 326392
rect 300584 326340 300636 326392
rect 300860 326340 300912 326392
rect 301688 326340 301740 326392
rect 321652 326340 321704 326392
rect 322480 326340 322532 326392
rect 322940 326340 322992 326392
rect 323584 326340 323636 326392
rect 327264 326340 327316 326392
rect 328000 326340 328052 326392
rect 328644 326340 328696 326392
rect 329472 326340 329524 326392
rect 329932 326340 329984 326392
rect 330576 326340 330628 326392
rect 350540 326340 350592 326392
rect 351368 326340 351420 326392
rect 354772 326340 354824 326392
rect 355324 326340 355376 326392
rect 356060 326340 356112 326392
rect 357164 326340 357216 326392
rect 364616 326340 364668 326392
rect 419540 326340 419592 326392
rect 385040 326272 385092 326324
rect 386052 326272 386104 326324
rect 386604 326272 386656 326324
rect 387524 326272 387576 326324
rect 405740 326272 405792 326324
rect 406844 326272 406896 326324
rect 295524 326204 295576 326256
rect 410064 326204 410116 326256
rect 410892 326204 410944 326256
rect 305276 326000 305328 326052
rect 306104 326000 306156 326052
rect 371424 325728 371476 325780
rect 372160 325728 372212 325780
rect 205640 325048 205692 325100
rect 298284 325048 298336 325100
rect 164240 324980 164292 325032
rect 276664 324980 276716 325032
rect 40040 324912 40092 324964
rect 247316 324912 247368 324964
rect 363788 324912 363840 324964
rect 416780 324912 416832 324964
rect 408500 324504 408552 324556
rect 409052 324504 409104 324556
rect 407212 324232 407264 324284
rect 407948 324232 408000 324284
rect 408592 323824 408644 323876
rect 409420 323824 409472 323876
rect 128360 323620 128412 323672
rect 274824 323620 274876 323672
rect 89720 323552 89772 323604
rect 262588 323552 262640 323604
rect 280160 323552 280212 323604
rect 280896 323552 280948 323604
rect 295432 323552 295484 323604
rect 295616 323552 295668 323604
rect 325792 323552 325844 323604
rect 325976 323552 326028 323604
rect 397736 323552 397788 323604
rect 525800 323552 525852 323604
rect 358912 323212 358964 323264
rect 359740 323212 359792 323264
rect 369860 323144 369912 323196
rect 370688 323144 370740 323196
rect 380900 322736 380952 322788
rect 382004 322736 382056 322788
rect 357624 322600 357676 322652
rect 358268 322600 358320 322652
rect 358820 322532 358872 322584
rect 359096 322532 359148 322584
rect 189080 322260 189132 322312
rect 291936 322260 291988 322312
rect 51080 322192 51132 322244
rect 250536 322192 250588 322244
rect 397644 322192 397696 322244
rect 529940 322192 529992 322244
rect 387892 322124 387944 322176
rect 388260 322124 388312 322176
rect 295340 322056 295392 322108
rect 296168 322056 296220 322108
rect 329840 321580 329892 321632
rect 330208 321580 330260 321632
rect 364892 320968 364944 321020
rect 420920 320968 420972 321020
rect 385316 320900 385368 320952
rect 487160 320900 487212 320952
rect 176660 320832 176712 320884
rect 289912 320832 289964 320884
rect 292580 320832 292632 320884
rect 292764 320832 292816 320884
rect 306380 320832 306432 320884
rect 306564 320832 306616 320884
rect 413192 320832 413244 320884
rect 576124 320832 576176 320884
rect 248420 320764 248472 320816
rect 248604 320764 248656 320816
rect 3424 320084 3476 320136
rect 232504 320084 232556 320136
rect 367376 319472 367428 319524
rect 427820 319472 427872 319524
rect 223580 319404 223632 319456
rect 303804 319404 303856 319456
rect 386696 319404 386748 319456
rect 489920 319404 489972 319456
rect 370320 318112 370372 318164
rect 438860 318112 438912 318164
rect 226340 318044 226392 318096
rect 305184 318044 305236 318096
rect 386604 318044 386656 318096
rect 494060 318044 494112 318096
rect 122840 316684 122892 316736
rect 271972 316684 272024 316736
rect 387800 316684 387852 316736
rect 498200 316684 498252 316736
rect 394700 315256 394752 315308
rect 518900 315256 518952 315308
rect 391940 313896 391992 313948
rect 512000 313896 512052 313948
rect 171140 312604 171192 312656
rect 286416 312604 286468 312656
rect 64880 312536 64932 312588
rect 254124 312536 254176 312588
rect 368756 312536 368808 312588
rect 434720 312536 434772 312588
rect 400864 311108 400916 311160
rect 532700 311108 532752 311160
rect 135260 309816 135312 309868
rect 276204 309816 276256 309868
rect 81440 309748 81492 309800
rect 259736 309748 259788 309800
rect 406016 309748 406068 309800
rect 554780 309748 554832 309800
rect 132500 308456 132552 308508
rect 274824 308456 274876 308508
rect 74540 308388 74592 308440
rect 258356 308388 258408 308440
rect 408592 308388 408644 308440
rect 564440 308388 564492 308440
rect 207020 307096 207072 307148
rect 294604 307096 294656 307148
rect 60740 307028 60792 307080
rect 253204 307028 253256 307080
rect 409880 307028 409932 307080
rect 568580 307028 568632 307080
rect 3332 306280 3384 306332
rect 383016 306280 383068 306332
rect 371516 305668 371568 305720
rect 441620 305668 441672 305720
rect 390836 305600 390888 305652
rect 505100 305600 505152 305652
rect 209780 304308 209832 304360
rect 297456 304308 297508 304360
rect 53840 304240 53892 304292
rect 251364 304240 251416 304292
rect 379612 304240 379664 304292
rect 470600 304240 470652 304292
rect 157340 302948 157392 303000
rect 283196 302948 283248 303000
rect 25504 302880 25556 302932
rect 241796 302880 241848 302932
rect 146300 301452 146352 301504
rect 280436 301452 280488 301504
rect 393504 301452 393556 301504
rect 513380 301452 513432 301504
rect 143540 300092 143592 300144
rect 279056 300092 279108 300144
rect 397552 300092 397604 300144
rect 527180 300092 527232 300144
rect 424324 299412 424376 299464
rect 580172 299412 580224 299464
rect 365904 298732 365956 298784
rect 423772 298732 423824 298784
rect 400312 297372 400364 297424
rect 536840 297372 536892 297424
rect 403072 295944 403124 295996
rect 547880 295944 547932 295996
rect 407304 294584 407356 294636
rect 557540 294584 557592 294636
rect 2872 293904 2924 293956
rect 10324 293904 10376 293956
rect 413284 293224 413336 293276
rect 572812 293224 572864 293276
rect 147680 291796 147732 291848
rect 280344 291796 280396 291848
rect 398932 291796 398984 291848
rect 531320 291796 531372 291848
rect 136640 290436 136692 290488
rect 277584 290436 277636 290488
rect 402980 290436 403032 290488
rect 545120 290436 545172 290488
rect 179420 289144 179472 289196
rect 287704 289144 287756 289196
rect 35900 289076 35952 289128
rect 244924 289076 244976 289128
rect 405924 289076 405976 289128
rect 556160 289076 556212 289128
rect 139400 287648 139452 287700
rect 273904 287648 273956 287700
rect 411444 287648 411496 287700
rect 571984 287648 572036 287700
rect 178040 286356 178092 286408
rect 289176 286356 289228 286408
rect 354956 286356 355008 286408
rect 387800 286356 387852 286408
rect 118700 286288 118752 286340
rect 269764 286288 269816 286340
rect 378416 286288 378468 286340
rect 465172 286288 465224 286340
rect 182180 284996 182232 285048
rect 286324 284996 286376 285048
rect 356336 284996 356388 285048
rect 394700 284996 394752 285048
rect 62120 284928 62172 284980
rect 254032 284928 254084 284980
rect 285680 284928 285732 284980
rect 323216 284928 323268 284980
rect 381084 284928 381136 284980
rect 473360 284928 473412 284980
rect 184940 283636 184992 283688
rect 291384 283636 291436 283688
rect 360476 283636 360528 283688
rect 408592 283636 408644 283688
rect 10324 283568 10376 283620
rect 236092 283568 236144 283620
rect 390744 283568 390796 283620
rect 506480 283568 506532 283620
rect 195980 282208 196032 282260
rect 295524 282208 295576 282260
rect 363144 282208 363196 282260
rect 415400 282208 415452 282260
rect 121460 282140 121512 282192
rect 271144 282140 271196 282192
rect 394884 282140 394936 282192
rect 520280 282140 520332 282192
rect 200120 280848 200172 280900
rect 295984 280848 296036 280900
rect 365812 280848 365864 280900
rect 426440 280848 426492 280900
rect 16580 280780 16632 280832
rect 239404 280780 239456 280832
rect 404544 280780 404596 280832
rect 552020 280780 552072 280832
rect 296720 279624 296772 279676
rect 322204 279624 322256 279676
rect 202880 279488 202932 279540
rect 296996 279488 297048 279540
rect 103520 279420 103572 279472
rect 264244 279420 264296 279472
rect 372804 279420 372856 279472
rect 448520 279420 448572 279472
rect 213920 278060 213972 278112
rect 300952 278060 301004 278112
rect 85580 277992 85632 278044
rect 261116 277992 261168 278044
rect 374276 277992 374328 278044
rect 451280 277992 451332 278044
rect 220820 276700 220872 276752
rect 302332 276700 302384 276752
rect 69020 276632 69072 276684
rect 255596 276632 255648 276684
rect 375564 276632 375616 276684
rect 455420 276632 455472 276684
rect 231860 275340 231912 275392
rect 306564 275340 306616 275392
rect 11704 275272 11756 275324
rect 234712 275272 234764 275324
rect 376944 275272 376996 275324
rect 458180 275272 458232 275324
rect 274824 274048 274876 274100
rect 319076 274048 319128 274100
rect 129740 273912 129792 273964
rect 274640 273912 274692 273964
rect 376852 273912 376904 273964
rect 462320 273912 462372 273964
rect 460204 273164 460256 273216
rect 580172 273164 580224 273216
rect 150440 272484 150492 272536
rect 280252 272484 280304 272536
rect 359096 272484 359148 272536
rect 402980 272484 403032 272536
rect 153200 271124 153252 271176
rect 281724 271124 281776 271176
rect 381544 271124 381596 271176
rect 469220 271124 469272 271176
rect 161480 269764 161532 269816
rect 284484 269764 284536 269816
rect 383844 269764 383896 269816
rect 481640 269764 481692 269816
rect 165620 268336 165672 268388
rect 285864 268336 285916 268388
rect 383752 268336 383804 268388
rect 484400 268336 484452 268388
rect 3240 267656 3292 267708
rect 231124 267656 231176 267708
rect 222200 266976 222252 267028
rect 303712 266976 303764 267028
rect 385224 266976 385276 267028
rect 488540 266976 488592 267028
rect 168472 265616 168524 265668
rect 287244 265616 287296 265668
rect 386420 265616 386472 265668
rect 491300 265616 491352 265668
rect 172520 264188 172572 264240
rect 287152 264188 287204 264240
rect 387984 264188 388036 264240
rect 495440 264188 495492 264240
rect 183560 262828 183612 262880
rect 291292 262828 291344 262880
rect 389180 262828 389232 262880
rect 498292 262828 498344 262880
rect 292580 261536 292632 261588
rect 324596 261536 324648 261588
rect 186320 261468 186372 261520
rect 292764 261468 292816 261520
rect 354864 261468 354916 261520
rect 389180 261468 389232 261520
rect 389364 261468 389416 261520
rect 502340 261468 502392 261520
rect 190460 260108 190512 260160
rect 292856 260108 292908 260160
rect 356244 260108 356296 260160
rect 391940 260108 391992 260160
rect 392124 260108 392176 260160
rect 509240 260108 509292 260160
rect 445024 259360 445076 259412
rect 580172 259360 580224 259412
rect 193312 258680 193364 258732
rect 294144 258680 294196 258732
rect 367284 258680 367336 258732
rect 432052 258680 432104 258732
rect 197360 257320 197412 257372
rect 295432 257320 295484 257372
rect 393412 257320 393464 257372
rect 516140 257320 516192 257372
rect 204260 256028 204312 256080
rect 298192 256028 298244 256080
rect 41420 255960 41472 256012
rect 247224 255960 247276 256012
rect 357624 255960 357676 256012
rect 398932 255960 398984 256012
rect 399024 255960 399076 256012
rect 534080 255960 534132 256012
rect 3332 255212 3384 255264
rect 17224 255212 17276 255264
rect 208400 254600 208452 254652
rect 298376 254600 298428 254652
rect 34520 254532 34572 254584
rect 245844 254532 245896 254584
rect 359004 254532 359056 254584
rect 400312 254532 400364 254584
rect 400404 254532 400456 254584
rect 538220 254532 538272 254584
rect 299480 253376 299532 253428
rect 320824 253376 320876 253428
rect 211160 253240 211212 253292
rect 299756 253240 299808 253292
rect 24124 253172 24176 253224
rect 240324 253172 240376 253224
rect 404452 253172 404504 253224
rect 547972 253172 548024 253224
rect 303620 252016 303672 252068
rect 328736 252016 328788 252068
rect 226432 251880 226484 251932
rect 303896 251880 303948 251932
rect 29000 251812 29052 251864
rect 243084 251812 243136 251864
rect 408684 251812 408736 251864
rect 563060 251812 563112 251864
rect 229100 250520 229152 250572
rect 305092 250520 305144 250572
rect 20720 250452 20772 250504
rect 241704 250452 241756 250504
rect 364984 250452 365036 250504
rect 409880 250452 409932 250504
rect 410156 250452 410208 250504
rect 565820 250452 565872 250504
rect 276204 249160 276256 249212
rect 318984 249160 319036 249212
rect 133880 249024 133932 249076
rect 276112 249024 276164 249076
rect 410064 249024 410116 249076
rect 569960 249024 570012 249076
rect 233240 247732 233292 247784
rect 306472 247732 306524 247784
rect 6920 247664 6972 247716
rect 233976 247664 234028 247716
rect 385132 247664 385184 247716
rect 485780 247664 485832 247716
rect 386512 246372 386564 246424
rect 140780 246304 140832 246356
rect 277492 246304 277544 246356
rect 353484 246304 353536 246356
rect 386420 246304 386472 246356
rect 492680 246304 492732 246356
rect 423036 245556 423088 245608
rect 580172 245556 580224 245608
rect 143632 244876 143684 244928
rect 278964 244876 279016 244928
rect 151820 243516 151872 243568
rect 281632 243516 281684 243568
rect 387892 243516 387944 243568
rect 496820 243516 496872 243568
rect 154580 242156 154632 242208
rect 283104 242156 283156 242208
rect 389272 242156 389324 242208
rect 499580 242156 499632 242208
rect 3240 241408 3292 241460
rect 232596 241408 232648 241460
rect 230480 240728 230532 240780
rect 305276 240728 305328 240780
rect 390652 240728 390704 240780
rect 503720 240728 503772 240780
rect 158720 239368 158772 239420
rect 283012 239368 283064 239420
rect 392032 239368 392084 239420
rect 510620 239368 510672 239420
rect 167000 238008 167052 238060
rect 285772 238008 285824 238060
rect 394792 238008 394844 238060
rect 517520 238008 517572 238060
rect 180800 236648 180852 236700
rect 290004 236648 290056 236700
rect 396264 236648 396316 236700
rect 521660 236648 521712 236700
rect 187700 235220 187752 235272
rect 292672 235220 292724 235272
rect 396172 235220 396224 235272
rect 524420 235220 524472 235272
rect 191840 233860 191892 233912
rect 294052 233860 294104 233912
rect 397460 233860 397512 233912
rect 528560 233860 528612 233912
rect 429844 233180 429896 233232
rect 579620 233180 579672 233232
rect 131120 232500 131172 232552
rect 274732 232500 274784 232552
rect 201592 231072 201644 231124
rect 296812 231072 296864 231124
rect 401784 231072 401836 231124
rect 539600 231072 539652 231124
rect 209872 229712 209924 229764
rect 299664 229712 299716 229764
rect 401692 229712 401744 229764
rect 542360 229712 542412 229764
rect 212540 228352 212592 228404
rect 299572 228352 299624 228404
rect 405832 228352 405884 228404
rect 553400 228352 553452 228404
rect 219440 226992 219492 227044
rect 302424 226992 302476 227044
rect 407212 226992 407264 227044
rect 560300 226992 560352 227044
rect 142160 225564 142212 225616
rect 278872 225564 278924 225616
rect 409972 225564 410024 225616
rect 567200 225564 567252 225616
rect 96620 224204 96672 224256
rect 265164 224204 265216 224256
rect 411352 224204 411404 224256
rect 574100 224204 574152 224256
rect 100760 222844 100812 222896
rect 265072 222844 265124 222896
rect 403624 222844 403676 222896
rect 540980 222844 541032 222896
rect 33140 221416 33192 221468
rect 244464 221416 244516 221468
rect 44180 220056 44232 220108
rect 248604 220056 248656 220108
rect 436744 219376 436796 219428
rect 580172 219376 580224 219428
rect 48320 218696 48372 218748
rect 249984 218696 250036 218748
rect 52460 217268 52512 217320
rect 249892 217268 249944 217320
rect 59360 215908 59412 215960
rect 251824 215908 251876 215960
rect 2780 214956 2832 215008
rect 4896 214956 4948 215008
rect 66260 214548 66312 214600
rect 255504 214548 255556 214600
rect 18604 213188 18656 213240
rect 238944 213188 238996 213240
rect 84200 211760 84252 211812
rect 261024 211760 261076 211812
rect 86960 210400 87012 210452
rect 260932 210400 260984 210452
rect 102140 209040 102192 209092
rect 266544 209040 266596 209092
rect 104900 207612 104952 207664
rect 266452 207612 266504 207664
rect 479524 206932 479576 206984
rect 580172 206932 580224 206984
rect 27620 206252 27672 206304
rect 242992 206252 243044 206304
rect 30380 204892 30432 204944
rect 244372 204892 244424 204944
rect 13176 203532 13228 203584
rect 237564 203532 237616 203584
rect 3332 202784 3384 202836
rect 18696 202784 18748 202836
rect 56600 202104 56652 202156
rect 252652 202104 252704 202156
rect 63500 200744 63552 200796
rect 254216 200744 254268 200796
rect 67640 199384 67692 199436
rect 255412 199384 255464 199436
rect 70400 197956 70452 198008
rect 256884 197956 256936 198008
rect 77300 196596 77352 196648
rect 258264 196596 258316 196648
rect 88340 195236 88392 195288
rect 262404 195236 262456 195288
rect 92480 193808 92532 193860
rect 262312 193808 262364 193860
rect 428464 193128 428516 193180
rect 580172 193128 580224 193180
rect 95240 192448 95292 192500
rect 263784 192448 263836 192500
rect 3148 188980 3200 189032
rect 11796 188980 11848 189032
rect 263784 180072 263836 180124
rect 316316 180072 316368 180124
rect 435364 179324 435416 179376
rect 580172 179324 580224 179376
rect 421564 166948 421616 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 229744 164160 229796 164212
rect 427084 153144 427136 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 21364 150356 21416 150408
rect 424324 139340 424376 139392
rect 580172 139340 580224 139392
rect 420184 126896 420236 126948
rect 579620 126896 579672 126948
rect 438124 113092 438176 113144
rect 580172 113092 580224 113144
rect 432604 100648 432656 100700
rect 579712 100648 579764 100700
rect 3516 97928 3568 97980
rect 22744 97928 22796 97980
rect 418804 86912 418856 86964
rect 579988 86912 580040 86964
rect 3516 85484 3568 85536
rect 13084 85484 13136 85536
rect 425704 73108 425756 73160
rect 580172 73108 580224 73160
rect 44272 72428 44324 72480
rect 248512 72428 248564 72480
rect 3516 71612 3568 71664
rect 7564 71612 7616 71664
rect 155960 71000 156012 71052
rect 282920 71000 282972 71052
rect 52552 64132 52604 64184
rect 251272 64132 251324 64184
rect 69112 61344 69164 61396
rect 255320 61344 255372 61396
rect 431224 60664 431276 60716
rect 579804 60664 579856 60716
rect 98000 59984 98052 60036
rect 265256 59984 265308 60036
rect 3056 59304 3108 59356
rect 10416 59304 10468 59356
rect 85672 55836 85724 55888
rect 260840 55836 260892 55888
rect 160192 54476 160244 54528
rect 284392 54476 284444 54528
rect 151912 53048 151964 53100
rect 281540 53048 281592 53100
rect 138020 51688 138072 51740
rect 277676 51688 277728 51740
rect 347964 51688 348016 51740
rect 365812 51688 365864 51740
rect 149060 50328 149112 50380
rect 280160 50328 280212 50380
rect 2780 48968 2832 49020
rect 234620 48968 234672 49020
rect 251272 48968 251324 49020
rect 312084 48968 312136 49020
rect 244372 47540 244424 47592
rect 310704 47540 310756 47592
rect 353392 47540 353444 47592
rect 385132 47540 385184 47592
rect 417424 46860 417476 46912
rect 580172 46860 580224 46912
rect 241704 46180 241756 46232
rect 309324 46180 309376 46232
rect 237564 44820 237616 44872
rect 307852 44820 307904 44872
rect 135352 43392 135404 43444
rect 276020 43392 276072 43444
rect 194600 42032 194652 42084
rect 294236 42032 294288 42084
rect 398840 42032 398892 42084
rect 531412 42032 531464 42084
rect 185032 40672 185084 40724
rect 291476 40672 291528 40724
rect 198740 39312 198792 39364
rect 295340 39312 295392 39364
rect 169760 37884 169812 37936
rect 287336 37884 287388 37936
rect 162860 36524 162912 36576
rect 284576 36524 284628 36576
rect 411260 36524 411312 36576
rect 571340 36524 571392 36576
rect 126980 35164 127032 35216
rect 273352 35164 273404 35216
rect 282920 35164 282972 35216
rect 307024 35164 307076 35216
rect 73160 33736 73212 33788
rect 256792 33736 256844 33788
rect 264980 33736 265032 33788
rect 316224 33736 316276 33788
rect 3516 33056 3568 33108
rect 8944 33056 8996 33108
rect 55220 32376 55272 32428
rect 251180 32376 251232 32428
rect 258264 32376 258316 32428
rect 314752 32376 314804 32428
rect 357532 32376 357584 32428
rect 397460 32376 397512 32428
rect 400220 32376 400272 32428
rect 535460 32376 535512 32428
rect 49700 31016 49752 31068
rect 249800 31016 249852 31068
rect 251180 31016 251232 31068
rect 311992 31016 312044 31068
rect 358912 31016 358964 31068
rect 404452 31016 404504 31068
rect 247224 29656 247276 29708
rect 310612 29656 310664 29708
rect 60832 29588 60884 29640
rect 252744 29588 252796 29640
rect 310704 29588 310756 29640
rect 330116 29588 330168 29640
rect 354772 29588 354824 29640
rect 390744 29588 390796 29640
rect 408500 29588 408552 29640
rect 564532 29588 564584 29640
rect 356152 28364 356204 28416
rect 393412 28364 393464 28416
rect 242992 28228 243044 28280
rect 309232 28228 309284 28280
rect 393320 28228 393372 28280
rect 514852 28228 514904 28280
rect 240324 26868 240376 26920
rect 309416 26868 309468 26920
rect 350632 26868 350684 26920
rect 375564 26868 375616 26920
rect 390560 26868 390612 26920
rect 506572 26868 506624 26920
rect 262312 25576 262364 25628
rect 316132 25576 316184 25628
rect 218060 25508 218112 25560
rect 298744 25508 298796 25560
rect 358084 25508 358136 25560
rect 372804 25508 372856 25560
rect 385040 25508 385092 25560
rect 490012 25508 490064 25560
rect 268016 24148 268068 24200
rect 317604 24148 317656 24200
rect 127072 24080 127124 24132
rect 273536 24080 273588 24132
rect 360384 24080 360436 24132
rect 407212 24080 407264 24132
rect 256792 22788 256844 22840
rect 313372 22788 313424 22840
rect 144920 22720 144972 22772
rect 278780 22720 278832 22772
rect 356060 22720 356112 22772
rect 396172 22720 396224 22772
rect 37280 21360 37332 21412
rect 245752 21360 245804 21412
rect 252560 21360 252612 21412
rect 312176 21360 312228 21412
rect 352104 21360 352156 21412
rect 382464 21360 382516 21412
rect 396080 21360 396132 21412
rect 523040 21360 523092 21412
rect 3424 20612 3476 20664
rect 414940 20612 414992 20664
rect 259736 19932 259788 19984
rect 302976 19932 303028 19984
rect 248512 18640 248564 18692
rect 310796 18640 310848 18692
rect 13820 18572 13872 18624
rect 238852 18572 238904 18624
rect 238944 18572 238996 18624
rect 301504 18572 301556 18624
rect 307760 18572 307812 18624
rect 330024 18572 330076 18624
rect 347872 18572 347924 18624
rect 368756 18572 368808 18624
rect 370504 18572 370556 18624
rect 412824 18572 412876 18624
rect 234620 17348 234672 17400
rect 306656 17348 306708 17400
rect 360292 17348 360344 17400
rect 405832 17348 405884 17400
rect 255320 17280 255372 17332
rect 313464 17280 313516 17332
rect 306472 17212 306524 17264
rect 328644 17212 328696 17264
rect 346584 17212 346636 17264
rect 360292 17212 360344 17264
rect 405740 17212 405792 17264
rect 556252 17212 556304 17264
rect 260656 15920 260708 15972
rect 291844 15920 291896 15972
rect 116400 15852 116452 15904
rect 270684 15852 270736 15904
rect 279056 15852 279108 15904
rect 319444 15852 319496 15904
rect 358820 15852 358872 15904
rect 402520 15852 402572 15904
rect 404360 15852 404412 15904
rect 550272 15852 550324 15904
rect 112352 14764 112404 14816
rect 269304 14764 269356 14816
rect 109040 14696 109092 14748
rect 267924 14696 267976 14748
rect 93860 14628 93912 14680
rect 263692 14628 263744 14680
rect 91560 14560 91612 14612
rect 262220 14560 262272 14612
rect 80888 14492 80940 14544
rect 259644 14492 259696 14544
rect 313832 14492 313884 14544
rect 331496 14492 331548 14544
rect 77392 14424 77444 14476
rect 258172 14424 258224 14476
rect 268108 14424 268160 14476
rect 313924 14424 313976 14476
rect 352012 14424 352064 14476
rect 381176 14424 381228 14476
rect 383660 14424 383712 14476
rect 482376 14424 482428 14476
rect 118792 13336 118844 13388
rect 270776 13336 270828 13388
rect 114744 13268 114796 13320
rect 270592 13268 270644 13320
rect 111616 13200 111668 13252
rect 269212 13200 269264 13252
rect 108120 13132 108172 13184
rect 267832 13132 267884 13184
rect 363052 13132 363104 13184
rect 415492 13132 415544 13184
rect 93952 13064 94004 13116
rect 263600 13064 263652 13116
rect 270776 13064 270828 13116
rect 317512 13064 317564 13116
rect 350540 13064 350592 13116
rect 377312 13064 377364 13116
rect 407120 13064 407172 13116
rect 559288 13064 559340 13116
rect 126980 11772 127032 11824
rect 128176 11772 128228 11824
rect 160100 11772 160152 11824
rect 161296 11772 161348 11824
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 216864 11772 216916 11824
rect 300860 11772 300912 11824
rect 349344 11772 349396 11824
rect 374276 11772 374328 11824
rect 8760 11704 8812 11756
rect 237472 11704 237524 11756
rect 271972 11704 272024 11756
rect 318892 11704 318944 11756
rect 373264 11704 373316 11756
rect 414296 11704 414348 11756
rect 422944 11704 422996 11756
rect 523132 11704 523184 11756
rect 226340 11636 226392 11688
rect 227536 11636 227588 11688
rect 372712 10820 372764 10872
rect 445760 10820 445812 10872
rect 372620 10752 372672 10804
rect 448612 10752 448664 10804
rect 374184 10684 374236 10736
rect 453304 10684 453356 10736
rect 375472 10616 375524 10668
rect 456892 10616 456944 10668
rect 376760 10548 376812 10600
rect 459928 10548 459980 10600
rect 378324 10480 378376 10532
rect 463976 10480 464028 10532
rect 173900 10412 173952 10464
rect 288532 10412 288584 10464
rect 378232 10412 378284 10464
rect 467472 10412 467524 10464
rect 83280 10344 83332 10396
rect 259460 10344 259512 10396
rect 345112 10344 345164 10396
rect 357532 10344 357584 10396
rect 380992 10344 381044 10396
rect 474096 10344 474148 10396
rect 79232 10276 79284 10328
rect 259552 10276 259604 10328
rect 261760 10276 261812 10328
rect 314844 10276 314896 10328
rect 349252 10276 349304 10328
rect 371516 10276 371568 10328
rect 382372 10276 382424 10328
rect 478144 10276 478196 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 249984 9120 250036 9172
rect 297364 9120 297416 9172
rect 254676 9052 254728 9104
rect 305736 9052 305788 9104
rect 76196 8984 76248 9036
rect 258080 8984 258132 9036
rect 349160 8984 349212 9036
rect 370596 8984 370648 9036
rect 72608 8916 72660 8968
rect 256700 8916 256752 8968
rect 317328 8916 317380 8968
rect 332784 8916 332836 8968
rect 353300 8916 353352 8968
rect 383568 8916 383620 8968
rect 387064 8916 387116 8968
rect 398840 8916 398892 8968
rect 412732 8916 412784 8968
rect 577412 8916 577464 8968
rect 377404 8236 377456 8288
rect 378876 8236 378928 8288
rect 237012 7624 237064 7676
rect 304264 7624 304316 7676
rect 310244 7624 310296 7676
rect 329932 7624 329984 7676
rect 347780 7624 347832 7676
rect 367008 7624 367060 7676
rect 176752 7556 176804 7608
rect 288624 7556 288676 7608
rect 290188 7556 290240 7608
rect 315304 7556 315356 7608
rect 351920 7556 351972 7608
rect 379980 7556 380032 7608
rect 380900 7556 380952 7608
rect 476948 7556 477000 7608
rect 3424 6808 3476 6860
rect 14464 6808 14516 6860
rect 367192 6468 367244 6520
rect 430856 6468 430908 6520
rect 368664 6400 368716 6452
rect 434444 6400 434496 6452
rect 369952 6332 370004 6384
rect 437940 6332 437992 6384
rect 281908 6264 281960 6316
rect 321744 6264 321796 6316
rect 371332 6264 371384 6316
rect 441528 6264 441580 6316
rect 234712 6196 234764 6248
rect 305644 6196 305696 6248
rect 345020 6196 345072 6248
rect 359924 6196 359976 6248
rect 371424 6196 371476 6248
rect 445024 6196 445076 6248
rect 12348 6128 12400 6180
rect 237748 6128 237800 6180
rect 242900 6128 242952 6180
rect 302884 6128 302936 6180
rect 346492 6128 346544 6180
rect 364616 6128 364668 6180
rect 412640 6128 412692 6180
rect 576308 6128 576360 6180
rect 366364 5516 366416 5568
rect 368204 5516 368256 5568
rect 303160 5176 303212 5228
rect 328552 5176 328604 5228
rect 299664 5108 299716 5160
rect 327356 5108 327408 5160
rect 296076 5040 296128 5092
rect 325792 5040 325844 5092
rect 288992 4972 289044 5024
rect 323032 4972 323084 5024
rect 285404 4904 285456 4956
rect 323124 4904 323176 4956
rect 278320 4836 278372 4888
rect 320364 4836 320416 4888
rect 351184 4836 351236 4888
rect 356336 4836 356388 4888
rect 218152 4768 218204 4820
rect 233884 4768 233936 4820
rect 246396 4768 246448 4820
rect 289084 4768 289136 4820
rect 292580 4768 292632 4820
rect 324504 4768 324556 4820
rect 354680 4768 354732 4820
rect 391848 4768 391900 4820
rect 401600 4768 401652 4820
rect 540796 4768 540848 4820
rect 382924 4496 382976 4548
rect 384764 4496 384816 4548
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 176660 4156 176712 4208
rect 177856 4156 177908 4208
rect 345664 4156 345716 4208
rect 352840 4156 352892 4208
rect 103336 4088 103388 4140
rect 266636 4088 266688 4140
rect 305552 4088 305604 4140
rect 328460 4088 328512 4140
rect 333888 4088 333940 4140
rect 336832 4088 336884 4140
rect 367100 4088 367152 4140
rect 429660 4088 429712 4140
rect 46664 4020 46716 4072
rect 248696 4020 248748 4072
rect 301964 4020 302016 4072
rect 327264 4020 327316 4072
rect 332692 4020 332744 4072
rect 337108 4020 337160 4072
rect 340880 4020 340932 4072
rect 346952 4020 347004 4072
rect 368480 4020 368532 4072
rect 433248 4020 433300 4072
rect 43076 3952 43128 4004
rect 247040 3952 247092 4004
rect 298468 3952 298520 4004
rect 327172 3952 327224 4004
rect 330392 3952 330444 4004
rect 336924 3952 336976 4004
rect 368572 3952 368624 4004
rect 436744 3952 436796 4004
rect 39580 3884 39632 3936
rect 247132 3884 247184 3936
rect 294880 3884 294932 3936
rect 325884 3884 325936 3936
rect 369860 3884 369912 3936
rect 440332 3884 440384 3936
rect 35992 3816 36044 3868
rect 245936 3816 245988 3868
rect 291384 3816 291436 3868
rect 324412 3816 324464 3868
rect 329012 3816 329064 3868
rect 334164 3816 334216 3868
rect 342628 3816 342680 3868
rect 349252 3816 349304 3868
rect 371240 3816 371292 3868
rect 443828 3816 443880 3868
rect 32404 3748 32456 3800
rect 244280 3748 244332 3800
rect 287796 3748 287848 3800
rect 322940 3748 322992 3800
rect 326804 3748 326856 3800
rect 335452 3748 335504 3800
rect 342352 3748 342404 3800
rect 348056 3748 348108 3800
rect 374184 3748 374236 3800
rect 450912 3748 450964 3800
rect 576124 3748 576176 3800
rect 578608 3748 578660 3800
rect 28908 3680 28960 3732
rect 243176 3680 243228 3732
rect 284300 3680 284352 3732
rect 321652 3680 321704 3732
rect 323308 3680 323360 3732
rect 334072 3680 334124 3732
rect 342536 3680 342588 3732
rect 350448 3680 350500 3732
rect 375380 3680 375432 3732
rect 458088 3680 458140 3732
rect 25320 3612 25372 3664
rect 241612 3612 241664 3664
rect 280712 3612 280764 3664
rect 321836 3612 321888 3664
rect 325608 3612 325660 3664
rect 335544 3612 335596 3664
rect 346400 3612 346452 3664
rect 362316 3612 362368 3664
rect 378140 3612 378192 3664
rect 465172 3612 465224 3664
rect 24216 3544 24268 3596
rect 241520 3544 241572 3596
rect 268016 3544 268068 3596
rect 268476 3544 268528 3596
rect 271880 3544 271932 3596
rect 272064 3544 272116 3596
rect 273628 3544 273680 3596
rect 318800 3544 318852 3596
rect 322112 3544 322164 3596
rect 329012 3544 329064 3596
rect 5264 3476 5316 3528
rect 6184 3476 6236 3528
rect 4068 3408 4120 3460
rect 10324 3476 10376 3528
rect 11152 3476 11204 3528
rect 15844 3476 15896 3528
rect 18236 3476 18288 3528
rect 24124 3476 24176 3528
rect 1676 3340 1728 3392
rect 11704 3340 11756 3392
rect 20628 3340 20680 3392
rect 240416 3476 240468 3528
rect 270040 3476 270092 3528
rect 317696 3476 317748 3528
rect 319720 3476 319772 3528
rect 332600 3544 332652 3596
rect 342444 3544 342496 3596
rect 351644 3544 351696 3596
rect 360200 3544 360252 3596
rect 408408 3544 408460 3596
rect 414112 3544 414164 3596
rect 581000 3544 581052 3596
rect 331588 3476 331640 3528
rect 333244 3476 333296 3528
rect 337476 3476 337528 3528
rect 338396 3476 338448 3528
rect 338672 3476 338724 3528
rect 339592 3476 339644 3528
rect 339684 3476 339736 3528
rect 340972 3476 341024 3528
rect 343640 3476 343692 3528
rect 354036 3476 354088 3528
rect 357440 3476 357492 3528
rect 358728 3476 358780 3528
rect 374000 3476 374052 3528
rect 375288 3476 375340 3528
rect 379520 3476 379572 3528
rect 472256 3476 472308 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 13544 3272 13596 3324
rect 18604 3272 18656 3324
rect 19432 3272 19484 3324
rect 240232 3408 240284 3460
rect 266544 3408 266596 3460
rect 316040 3408 316092 3460
rect 318524 3408 318576 3460
rect 332784 3408 332836 3460
rect 343732 3408 343784 3460
rect 355232 3408 355284 3460
rect 361580 3408 361632 3460
rect 411904 3408 411956 3460
rect 415400 3408 415452 3460
rect 416688 3408 416740 3460
rect 416780 3408 416832 3460
rect 582196 3408 582248 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 77300 3340 77352 3392
rect 78220 3340 78272 3392
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 106924 3340 106976 3392
rect 268200 3340 268252 3392
rect 309048 3340 309100 3392
rect 329840 3340 329892 3392
rect 341064 3340 341116 3392
rect 344560 3340 344612 3392
rect 365720 3340 365772 3392
rect 426164 3340 426216 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 118700 3272 118752 3324
rect 119896 3272 119948 3324
rect 9956 3204 10008 3256
rect 13176 3204 13228 3256
rect 114008 3204 114060 3256
rect 269120 3272 269172 3324
rect 312636 3272 312688 3324
rect 331404 3272 331456 3324
rect 364432 3272 364484 3324
rect 422576 3272 422628 3324
rect 121092 3204 121144 3256
rect 271880 3204 271932 3256
rect 315028 3204 315080 3256
rect 331220 3204 331272 3256
rect 364340 3204 364392 3256
rect 418988 3204 419040 3256
rect 23020 3136 23072 3188
rect 25504 3136 25556 3188
rect 218060 3136 218112 3188
rect 219256 3136 219308 3188
rect 234620 3136 234672 3188
rect 235816 3136 235868 3188
rect 316224 3136 316276 3188
rect 331312 3136 331364 3188
rect 336280 3136 336332 3188
rect 338212 3136 338264 3188
rect 398932 3136 398984 3188
rect 400128 3136 400180 3188
rect 414020 3136 414072 3188
rect 416780 3136 416832 3188
rect 572 3068 624 3120
rect 4804 3068 4856 3120
rect 329196 3000 329248 3052
rect 335636 3000 335688 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 341156 2864 341208 2916
rect 345756 2864 345808 2916
rect 299480 2048 299532 2100
rect 300768 2048 300820 2100
rect 423680 960 423732 1012
rect 424968 960 425020 1012
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3344 618322 3372 619103
rect 3332 618316 3384 618322
rect 3332 618258 3384 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3436 460193 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3528 465746 3556 632023
rect 3606 580000 3662 580009
rect 3606 579935 3662 579944
rect 3620 465882 3648 579935
rect 3698 527912 3754 527921
rect 3698 527847 3754 527856
rect 3712 466018 3740 527847
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3712 465990 3832 466018
rect 3620 465854 3740 465882
rect 3528 465718 3648 465746
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3620 460426 3648 465718
rect 3608 460420 3660 460426
rect 3608 460362 3660 460368
rect 3712 460358 3740 465854
rect 3700 460352 3752 460358
rect 3700 460294 3752 460300
rect 3804 460290 3832 465990
rect 3792 460284 3844 460290
rect 3792 460226 3844 460232
rect 3896 460222 3924 475623
rect 4896 460964 4948 460970
rect 4896 460906 4948 460912
rect 3884 460216 3936 460222
rect 3422 460184 3478 460193
rect 3884 460158 3936 460164
rect 3422 460119 3478 460128
rect 3516 458244 3568 458250
rect 3516 458186 3568 458192
rect 3424 457496 3476 457502
rect 3424 457438 3476 457444
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3436 397497 3464 457438
rect 3528 423609 3556 458186
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3514 337376 3570 337385
rect 3514 337311 3570 337320
rect 3424 320136 3476 320142
rect 3424 320078 3476 320084
rect 3436 319297 3464 320078
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3422 313984 3478 313993
rect 3422 313919 3478 313928
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2872 293956 2924 293962
rect 2872 293898 2924 293904
rect 2884 293185 2912 293898
rect 2870 293176 2926 293185
rect 2870 293111 2926 293120
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3332 255264 3384 255270
rect 3332 255206 3384 255212
rect 3344 254153 3372 255206
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 2780 215008 2832 215014
rect 2778 214976 2780 214985
rect 2832 214976 2834 214985
rect 2778 214911 2834 214920
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2780 49020 2832 49026
rect 2780 48962 2832 48968
rect 2792 16574 2820 48962
rect 3436 45529 3464 313919
rect 3528 110673 3556 337311
rect 4804 326392 4856 326398
rect 4804 326334 4856 326340
rect 3606 316704 3662 316713
rect 3606 316639 3662 316648
rect 3620 136785 3648 316639
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 3514 110664 3570 110673
rect 3514 110599 3570 110608
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2792 16546 2912 16574
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 572 3120 624 3126
rect 572 3062 624 3068
rect 584 480 612 3062
rect 1688 480 1716 3334
rect 2884 480 2912 16546
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 4816 3126 4844 326334
rect 4908 215014 4936 460906
rect 40052 460329 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 104912 468518 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 104900 468512 104952 468518
rect 104900 468454 104952 468460
rect 136652 460630 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700602 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700596 154172 700602
rect 154120 700538 154172 700544
rect 169772 467158 169800 702406
rect 169760 467152 169812 467158
rect 169760 467094 169812 467100
rect 201512 460834 201540 702986
rect 218992 700670 219020 703520
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 235184 698970 235212 703520
rect 235172 698964 235224 698970
rect 235172 698906 235224 698912
rect 267660 697610 267688 703520
rect 283852 700806 283880 703520
rect 283840 700800 283892 700806
rect 283840 700742 283892 700748
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 226984 462528 227036 462534
rect 226984 462470 227036 462476
rect 225604 462460 225656 462466
rect 225604 462402 225656 462408
rect 201500 460828 201552 460834
rect 201500 460770 201552 460776
rect 136640 460624 136692 460630
rect 136640 460566 136692 460572
rect 40038 460320 40094 460329
rect 40038 460255 40094 460264
rect 225616 358766 225644 462402
rect 226996 411262 227024 462470
rect 233976 461372 234028 461378
rect 233976 461314 234028 461320
rect 228364 461100 228416 461106
rect 228364 461042 228416 461048
rect 226984 411256 227036 411262
rect 226984 411198 227036 411204
rect 225604 358760 225656 358766
rect 225604 358702 225656 358708
rect 228376 346390 228404 461042
rect 229744 461032 229796 461038
rect 229744 460974 229796 460980
rect 228364 346384 228416 346390
rect 228364 346326 228416 346332
rect 124220 336388 124272 336394
rect 124220 336330 124272 336336
rect 117320 336320 117372 336326
rect 117320 336262 117372 336268
rect 110420 336252 110472 336258
rect 110420 336194 110472 336200
rect 99380 336184 99432 336190
rect 99380 336126 99432 336132
rect 15844 336116 15896 336122
rect 15844 336058 15896 336064
rect 6184 336048 6236 336054
rect 6184 335990 6236 335996
rect 4896 215008 4948 215014
rect 4896 214950 4948 214956
rect 6196 3534 6224 335990
rect 7562 334656 7618 334665
rect 7562 334591 7618 334600
rect 6920 247716 6972 247722
rect 6920 247658 6972 247664
rect 6932 16574 6960 247658
rect 7576 71670 7604 334591
rect 8942 333296 8998 333305
rect 8942 333231 8998 333240
rect 7564 71664 7616 71670
rect 7564 71606 7616 71612
rect 8956 33114 8984 333231
rect 10322 320784 10378 320793
rect 10322 320719 10378 320728
rect 10336 293962 10364 320719
rect 11794 318064 11850 318073
rect 11794 317999 11850 318008
rect 10324 293956 10376 293962
rect 10324 293898 10376 293904
rect 10414 293176 10470 293185
rect 10414 293111 10470 293120
rect 10324 283620 10376 283626
rect 10324 283562 10376 283568
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 6932 16546 7696 16574
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 5276 480 5304 3470
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 16546
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 480 8800 11698
rect 10336 3534 10364 283562
rect 10428 59362 10456 293111
rect 11704 275324 11756 275330
rect 11704 275266 11756 275272
rect 10416 59356 10468 59362
rect 10416 59298 10468 59304
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 9956 3256 10008 3262
rect 9956 3198 10008 3204
rect 9968 480 9996 3198
rect 11164 480 11192 3470
rect 11716 3398 11744 275266
rect 11808 189038 11836 317999
rect 13082 315344 13138 315353
rect 13082 315279 13138 315288
rect 11796 189032 11848 189038
rect 11796 188974 11848 188980
rect 13096 85542 13124 315279
rect 14462 311128 14518 311137
rect 14462 311063 14518 311072
rect 13176 203584 13228 203590
rect 13176 203526 13228 203532
rect 13084 85536 13136 85542
rect 13084 85478 13136 85484
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 12360 480 12388 6122
rect 13188 3262 13216 203526
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13832 16574 13860 18566
rect 13832 16546 14320 16574
rect 13544 3324 13596 3330
rect 13544 3266 13596 3272
rect 13176 3256 13228 3262
rect 13176 3198 13228 3204
rect 13556 480 13584 3266
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 6866 14504 311063
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 15856 3534 15884 336058
rect 46940 331900 46992 331906
rect 46940 331842 46992 331848
rect 26240 329112 26292 329118
rect 26240 329054 26292 329060
rect 25504 302932 25556 302938
rect 25504 302874 25556 302880
rect 17222 298752 17278 298761
rect 17222 298687 17278 298696
rect 16580 280832 16632 280838
rect 16580 280774 16632 280780
rect 16592 16574 16620 280774
rect 17236 255270 17264 298687
rect 18694 297392 18750 297401
rect 18694 297327 18750 297336
rect 17224 255264 17276 255270
rect 17224 255206 17276 255212
rect 18604 213240 18656 213246
rect 18604 213182 18656 213188
rect 16592 16546 17080 16574
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15934 3496 15990 3505
rect 15934 3431 15990 3440
rect 15948 480 15976 3431
rect 17052 480 17080 16546
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 480 18276 3470
rect 18616 3330 18644 213182
rect 18708 202842 18736 297327
rect 21362 296032 21418 296041
rect 21362 295967 21418 295976
rect 20720 250504 20772 250510
rect 20720 250446 20772 250452
rect 18696 202836 18748 202842
rect 18696 202778 18748 202784
rect 20732 16574 20760 250446
rect 21376 150414 21404 295967
rect 22742 294536 22798 294545
rect 22742 294471 22798 294480
rect 21364 150408 21416 150414
rect 21364 150350 21416 150356
rect 22756 97986 22784 294471
rect 24124 253224 24176 253230
rect 24124 253166 24176 253172
rect 22744 97980 22796 97986
rect 22744 97922 22796 97928
rect 20732 16546 21864 16574
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 18604 3324 18656 3330
rect 18604 3266 18656 3272
rect 19432 3324 19484 3330
rect 19432 3266 19484 3272
rect 19444 480 19472 3266
rect 20640 480 20668 3334
rect 21836 480 21864 16546
rect 24136 3534 24164 253166
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23032 480 23060 3130
rect 24228 480 24256 3538
rect 25332 480 25360 3606
rect 25516 3194 25544 302874
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 329054
rect 40040 324964 40092 324970
rect 40040 324906 40092 324912
rect 35900 289128 35952 289134
rect 35900 289070 35952 289076
rect 34520 254584 34572 254590
rect 34520 254526 34572 254532
rect 29000 251864 29052 251870
rect 29000 251806 29052 251812
rect 27620 206304 27672 206310
rect 27620 206246 27672 206252
rect 27632 16574 27660 206246
rect 29012 16574 29040 251806
rect 33140 221468 33192 221474
rect 33140 221410 33192 221416
rect 30380 204944 30432 204950
rect 30380 204886 30432 204892
rect 30392 16574 30420 204886
rect 33152 16574 33180 221410
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 28920 480 28948 3674
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32416 480 32444 3742
rect 33612 480 33640 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 254526
rect 35912 16574 35940 289070
rect 37280 21412 37332 21418
rect 37280 21354 37332 21360
rect 37292 16574 37320 21354
rect 40052 16574 40080 324906
rect 41420 256012 41472 256018
rect 41420 255954 41472 255960
rect 41432 16574 41460 255954
rect 44180 220108 44232 220114
rect 44180 220050 44232 220056
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35992 3868 36044 3874
rect 35992 3810 36044 3816
rect 36004 480 36032 3810
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39592 480 39620 3878
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 44192 6914 44220 220050
rect 44272 72480 44324 72486
rect 44272 72422 44324 72428
rect 44284 16574 44312 72422
rect 46952 16574 46980 331842
rect 57980 330540 58032 330546
rect 57980 330482 58032 330488
rect 51080 322244 51132 322250
rect 51080 322186 51132 322192
rect 48320 218748 48372 218754
rect 48320 218690 48372 218696
rect 48332 16574 48360 218690
rect 49700 31068 49752 31074
rect 49700 31010 49752 31016
rect 49712 16574 49740 31010
rect 44284 16546 45048 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 43076 4004 43128 4010
rect 43076 3946 43128 3952
rect 43088 480 43116 3946
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 46676 480 46704 4014
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 322186
rect 53840 304292 53892 304298
rect 53840 304234 53892 304240
rect 52460 217320 52512 217326
rect 52460 217262 52512 217268
rect 52472 6914 52500 217262
rect 52552 64184 52604 64190
rect 52552 64126 52604 64132
rect 52564 16574 52592 64126
rect 53852 16574 53880 304234
rect 56600 202156 56652 202162
rect 56600 202098 56652 202104
rect 55220 32428 55272 32434
rect 55220 32370 55272 32376
rect 55232 16574 55260 32370
rect 56612 16574 56640 202098
rect 57992 16574 58020 330482
rect 89720 323604 89772 323610
rect 89720 323546 89772 323552
rect 64880 312588 64932 312594
rect 64880 312530 64932 312536
rect 60740 307080 60792 307086
rect 60740 307022 60792 307028
rect 59360 215960 59412 215966
rect 59360 215902 59412 215908
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 215902
rect 60752 3398 60780 307022
rect 62120 284980 62172 284986
rect 62120 284922 62172 284928
rect 60832 29640 60884 29646
rect 60832 29582 60884 29588
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 29582
rect 62132 16574 62160 284922
rect 63500 200796 63552 200802
rect 63500 200738 63552 200744
rect 63512 16574 63540 200738
rect 64892 16574 64920 312530
rect 81440 309800 81492 309806
rect 81440 309742 81492 309748
rect 74540 308440 74592 308446
rect 74540 308382 74592 308388
rect 69020 276684 69072 276690
rect 69020 276626 69072 276632
rect 66260 214600 66312 214606
rect 66260 214542 66312 214548
rect 66272 16574 66300 214542
rect 67640 199436 67692 199442
rect 67640 199378 67692 199384
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 199378
rect 69032 6914 69060 276626
rect 70400 198008 70452 198014
rect 70400 197950 70452 197956
rect 69112 61396 69164 61402
rect 69112 61338 69164 61344
rect 69124 16574 69152 61338
rect 70412 16574 70440 197950
rect 73160 33788 73212 33794
rect 73160 33730 73212 33736
rect 73172 16574 73200 33730
rect 74552 16574 74580 308382
rect 77300 196648 77352 196654
rect 77300 196590 77352 196596
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72608 8968 72660 8974
rect 72608 8910 72660 8916
rect 72620 480 72648 8910
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 76196 9036 76248 9042
rect 76196 8978 76248 8984
rect 76208 480 76236 8978
rect 77312 3398 77340 196590
rect 81452 16574 81480 309742
rect 85580 278044 85632 278050
rect 85580 277986 85632 277992
rect 84200 211812 84252 211818
rect 84200 211754 84252 211760
rect 81452 16546 81664 16574
rect 80888 14544 80940 14550
rect 80888 14486 80940 14492
rect 77392 14476 77444 14482
rect 77392 14418 77444 14424
rect 77300 3392 77352 3398
rect 77300 3334 77352 3340
rect 77404 480 77432 14418
rect 79232 10328 79284 10334
rect 79232 10270 79284 10276
rect 78220 3392 78272 3398
rect 78220 3334 78272 3340
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78232 354 78260 3334
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 10270
rect 80900 480 80928 14486
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 10396 83332 10402
rect 83280 10338 83332 10344
rect 83292 480 83320 10338
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 211754
rect 85592 3398 85620 277986
rect 86960 210452 87012 210458
rect 86960 210394 87012 210400
rect 85672 55888 85724 55894
rect 85672 55830 85724 55836
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 85684 480 85712 55830
rect 86972 16574 87000 210394
rect 88340 195288 88392 195294
rect 88340 195230 88392 195236
rect 88352 16574 88380 195230
rect 89732 16574 89760 323546
rect 96620 224256 96672 224262
rect 96620 224198 96672 224204
rect 92480 193860 92532 193866
rect 92480 193802 92532 193808
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 14612 91612 14618
rect 91560 14554 91612 14560
rect 91572 480 91600 14554
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 193802
rect 95240 192500 95292 192506
rect 95240 192442 95292 192448
rect 95252 16574 95280 192442
rect 96632 16574 96660 224198
rect 98000 60036 98052 60042
rect 98000 59978 98052 59984
rect 98012 16574 98040 59978
rect 99392 16574 99420 336126
rect 103520 279472 103572 279478
rect 103520 279414 103572 279420
rect 100760 222896 100812 222902
rect 100760 222838 100812 222844
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93860 14680 93912 14686
rect 93860 14622 93912 14628
rect 93872 3398 93900 14622
rect 93952 13116 94004 13122
rect 93952 13058 94004 13064
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 13058
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 222838
rect 102140 209092 102192 209098
rect 102140 209034 102192 209040
rect 102152 16574 102180 209034
rect 103532 16574 103560 279414
rect 104900 207664 104952 207670
rect 104900 207606 104952 207612
rect 104912 16574 104940 207606
rect 110432 16574 110460 336194
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 110432 16546 110552 16574
rect 102244 480 102272 16546
rect 103336 4140 103388 4146
rect 103336 4082 103388 4088
rect 103348 480 103376 4082
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 109040 14748 109092 14754
rect 109040 14690 109092 14696
rect 108120 13184 108172 13190
rect 108120 13126 108172 13132
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 106936 480 106964 3334
rect 108132 480 108160 13126
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 14690
rect 110524 480 110552 16546
rect 116400 15904 116452 15910
rect 116400 15846 116452 15852
rect 112352 14816 112404 14822
rect 112352 14758 112404 14764
rect 111616 13252 111668 13258
rect 111616 13194 111668 13200
rect 111628 480 111656 13194
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 14758
rect 114744 13320 114796 13326
rect 114744 13262 114796 13268
rect 114008 3256 114060 3262
rect 114008 3198 114060 3204
rect 114020 480 114048 3198
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 13262
rect 116412 480 116440 15846
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 336262
rect 122840 316736 122892 316742
rect 122840 316678 122892 316684
rect 118700 286340 118752 286346
rect 118700 286282 118752 286288
rect 118712 3330 118740 286282
rect 121460 282192 121512 282198
rect 121460 282134 121512 282140
rect 121472 16574 121500 282134
rect 122852 16574 122880 316678
rect 124232 16574 124260 336330
rect 224960 334620 225012 334626
rect 224960 334562 225012 334568
rect 175280 331968 175332 331974
rect 175280 331910 175332 331916
rect 168380 330608 168432 330614
rect 168380 330550 168432 330556
rect 160100 329180 160152 329186
rect 160100 329122 160152 329128
rect 125600 327752 125652 327758
rect 125600 327694 125652 327700
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118792 13388 118844 13394
rect 118792 13330 118844 13336
rect 118700 3324 118752 3330
rect 118700 3266 118752 3272
rect 118804 480 118832 13330
rect 119896 3324 119948 3330
rect 119896 3266 119948 3272
rect 119908 480 119936 3266
rect 121092 3256 121144 3262
rect 121092 3198 121144 3204
rect 121104 480 121132 3198
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 327694
rect 128360 323672 128412 323678
rect 128360 323614 128412 323620
rect 126980 35216 127032 35222
rect 126980 35158 127032 35164
rect 126992 11830 127020 35158
rect 127072 24132 127124 24138
rect 127072 24074 127124 24080
rect 126980 11824 127032 11830
rect 126980 11766 127032 11772
rect 127084 6914 127112 24074
rect 128372 16574 128400 323614
rect 135260 309868 135312 309874
rect 135260 309810 135312 309816
rect 132500 308508 132552 308514
rect 132500 308450 132552 308456
rect 129740 273964 129792 273970
rect 129740 273906 129792 273912
rect 129752 16574 129780 273906
rect 131120 232552 131172 232558
rect 131120 232494 131172 232500
rect 131132 16574 131160 232494
rect 132512 16574 132540 308450
rect 133880 249076 133932 249082
rect 133880 249018 133932 249024
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128176 11824 128228 11830
rect 128176 11766 128228 11772
rect 126992 6886 127112 6914
rect 126992 480 127020 6886
rect 128188 480 128216 11766
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 249018
rect 135272 4214 135300 309810
rect 157340 303000 157392 303006
rect 157340 302942 157392 302948
rect 146300 301504 146352 301510
rect 146300 301446 146352 301452
rect 143540 300144 143592 300150
rect 143540 300086 143592 300092
rect 136640 290488 136692 290494
rect 136640 290430 136692 290436
rect 135352 43444 135404 43450
rect 135352 43386 135404 43392
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 135364 3482 135392 43386
rect 136652 16574 136680 290430
rect 139400 287700 139452 287706
rect 139400 287642 139452 287648
rect 138020 51740 138072 51746
rect 138020 51682 138072 51688
rect 138032 16574 138060 51682
rect 139412 16574 139440 287642
rect 140780 246356 140832 246362
rect 140780 246298 140832 246304
rect 140792 16574 140820 246298
rect 142160 225616 142212 225622
rect 142160 225558 142212 225564
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 4150
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 225558
rect 143552 480 143580 300086
rect 143632 244928 143684 244934
rect 143632 244870 143684 244876
rect 143644 16574 143672 244870
rect 144920 22772 144972 22778
rect 144920 22714 144972 22720
rect 144932 16574 144960 22714
rect 146312 16574 146340 301446
rect 147680 291848 147732 291854
rect 147680 291790 147732 291796
rect 147692 16574 147720 291790
rect 150440 272536 150492 272542
rect 150440 272478 150492 272484
rect 149060 50380 149112 50386
rect 149060 50322 149112 50328
rect 149072 16574 149100 50322
rect 150452 16574 150480 272478
rect 153200 271176 153252 271182
rect 153200 271118 153252 271124
rect 151820 243568 151872 243574
rect 151820 243510 151872 243516
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 243510
rect 151912 53100 151964 53106
rect 151912 53042 151964 53048
rect 151924 16574 151952 53042
rect 153212 16574 153240 271118
rect 154580 242208 154632 242214
rect 154580 242150 154632 242156
rect 154592 16574 154620 242150
rect 155960 71052 156012 71058
rect 155960 70994 156012 71000
rect 155972 16574 156000 70994
rect 157352 16574 157380 302942
rect 158720 239420 158772 239426
rect 158720 239362 158772 239368
rect 158732 16574 158760 239362
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11830 160140 329122
rect 164240 325032 164292 325038
rect 164240 324974 164292 324980
rect 161480 269816 161532 269822
rect 161480 269758 161532 269764
rect 160192 54528 160244 54534
rect 160192 54470 160244 54476
rect 160100 11824 160152 11830
rect 160100 11766 160152 11772
rect 160204 6914 160232 54470
rect 161492 16574 161520 269758
rect 162860 36576 162912 36582
rect 162860 36518 162912 36524
rect 162872 16574 162900 36518
rect 164252 16574 164280 324974
rect 165620 268388 165672 268394
rect 165620 268330 165672 268336
rect 165632 16574 165660 268330
rect 167000 238060 167052 238066
rect 167000 238002 167052 238008
rect 167012 16574 167040 238002
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11824 161348 11830
rect 161296 11766 161348 11772
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11766
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 330550
rect 171140 312656 171192 312662
rect 171140 312598 171192 312604
rect 168472 265668 168524 265674
rect 168472 265610 168524 265616
rect 168484 16574 168512 265610
rect 169760 37936 169812 37942
rect 169760 37878 169812 37884
rect 169772 16574 169800 37878
rect 171152 16574 171180 312598
rect 172520 264240 172572 264246
rect 172520 264182 172572 264188
rect 172532 16574 172560 264182
rect 175292 16574 175320 331910
rect 201500 329248 201552 329254
rect 201500 329190 201552 329196
rect 193220 326460 193272 326466
rect 193220 326402 193272 326408
rect 189080 322312 189132 322318
rect 189080 322254 189132 322260
rect 176660 320884 176712 320890
rect 176660 320826 176712 320832
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 175292 16546 175504 16574
rect 169588 480 169616 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173900 10464 173952 10470
rect 173900 10406 173952 10412
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 10406
rect 175476 480 175504 16546
rect 176672 4214 176700 320826
rect 179420 289196 179472 289202
rect 179420 289138 179472 289144
rect 178040 286408 178092 286414
rect 178040 286350 178092 286356
rect 178052 16574 178080 286350
rect 179432 16574 179460 289138
rect 182180 285048 182232 285054
rect 182180 284990 182232 284996
rect 180800 236700 180852 236706
rect 180800 236642 180852 236648
rect 180812 16574 180840 236642
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 176752 7608 176804 7614
rect 176752 7550 176804 7556
rect 176660 4208 176712 4214
rect 176660 4150 176712 4156
rect 176764 3482 176792 7550
rect 177856 4208 177908 4214
rect 177856 4150 177908 4156
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 4150
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 284990
rect 184940 283688 184992 283694
rect 184940 283630 184992 283636
rect 183560 262880 183612 262886
rect 183560 262822 183612 262828
rect 183572 16574 183600 262822
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 283630
rect 186320 261520 186372 261526
rect 186320 261462 186372 261468
rect 185032 40724 185084 40730
rect 185032 40666 185084 40672
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 185044 6914 185072 40666
rect 186332 16574 186360 261462
rect 187700 235272 187752 235278
rect 187700 235214 187752 235220
rect 187712 16574 187740 235214
rect 189092 16574 189120 322254
rect 190460 260160 190512 260166
rect 190460 260102 190512 260108
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 260102
rect 191840 233912 191892 233918
rect 191840 233854 191892 233860
rect 191852 16574 191880 233854
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 326402
rect 195980 282260 196032 282266
rect 195980 282202 196032 282208
rect 193312 258732 193364 258738
rect 193312 258674 193364 258680
rect 193324 16574 193352 258674
rect 194600 42084 194652 42090
rect 194600 42026 194652 42032
rect 194612 16574 194640 42026
rect 195992 16574 196020 282202
rect 200120 280900 200172 280906
rect 200120 280842 200172 280848
rect 197360 257372 197412 257378
rect 197360 257314 197412 257320
rect 197372 16574 197400 257314
rect 198740 39364 198792 39370
rect 198740 39306 198792 39312
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 39306
rect 200132 16574 200160 280842
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 329190
rect 215300 327820 215352 327826
rect 215300 327762 215352 327768
rect 205640 325100 205692 325106
rect 205640 325042 205692 325048
rect 202880 279540 202932 279546
rect 202880 279482 202932 279488
rect 201592 231124 201644 231130
rect 201592 231066 201644 231072
rect 201604 16574 201632 231066
rect 202892 16574 202920 279482
rect 204260 256080 204312 256086
rect 204260 256022 204312 256028
rect 204272 16574 204300 256022
rect 205652 16574 205680 325042
rect 207020 307148 207072 307154
rect 207020 307090 207072 307096
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 307090
rect 209780 304360 209832 304366
rect 209780 304302 209832 304308
rect 208400 254652 208452 254658
rect 208400 254594 208452 254600
rect 208412 16574 208440 254594
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 304302
rect 213920 278112 213972 278118
rect 213920 278054 213972 278060
rect 211160 253292 211212 253298
rect 211160 253234 211212 253240
rect 209872 229764 209924 229770
rect 209872 229706 209924 229712
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 229706
rect 211172 16574 211200 253234
rect 212540 228404 212592 228410
rect 212540 228346 212592 228352
rect 212552 16574 212580 228346
rect 213932 16574 213960 278054
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 327762
rect 223580 319456 223632 319462
rect 223580 319398 223632 319404
rect 220820 276752 220872 276758
rect 220820 276694 220872 276700
rect 219440 227044 219492 227050
rect 219440 226986 219492 226992
rect 218060 25560 218112 25566
rect 218060 25502 218112 25508
rect 216864 11824 216916 11830
rect 216864 11766 216916 11772
rect 216876 480 216904 11766
rect 218072 3194 218100 25502
rect 219452 16574 219480 226986
rect 220832 16574 220860 276694
rect 222200 267028 222252 267034
rect 222200 266970 222252 266976
rect 222212 16574 222240 266970
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 218152 4820 218204 4826
rect 218152 4762 218204 4768
rect 218060 3188 218112 3194
rect 218060 3130 218112 3136
rect 218164 2394 218192 4762
rect 219256 3188 219308 3194
rect 219256 3130 219308 3136
rect 218072 2366 218192 2394
rect 218072 480 218100 2366
rect 219268 480 219296 3130
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 319398
rect 224972 16574 225000 334562
rect 227720 333260 227772 333266
rect 227720 333202 227772 333208
rect 226340 318096 226392 318102
rect 226340 318038 226392 318044
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 11694 226380 318038
rect 226432 251932 226484 251938
rect 226432 251874 226484 251880
rect 226340 11688 226392 11694
rect 226340 11630 226392 11636
rect 226444 6914 226472 251874
rect 227732 16574 227760 333202
rect 229100 250572 229152 250578
rect 229100 250514 229152 250520
rect 229112 16574 229140 250514
rect 229756 164218 229784 460974
rect 233884 458856 233936 458862
rect 233884 458798 233936 458804
rect 232504 458652 232556 458658
rect 232504 458594 232556 458600
rect 231124 458584 231176 458590
rect 231124 458526 231176 458532
rect 231136 267714 231164 458526
rect 232516 320142 232544 458594
rect 233896 372570 233924 458798
rect 233988 449886 234016 461314
rect 266372 460154 266400 697546
rect 298100 643136 298152 643142
rect 298100 643078 298152 643084
rect 296720 616888 296772 616894
rect 296720 616830 296772 616836
rect 293960 590708 294012 590714
rect 293960 590650 294012 590656
rect 292580 563100 292632 563106
rect 292580 563042 292632 563048
rect 288440 536852 288492 536858
rect 288440 536794 288492 536800
rect 287060 510672 287112 510678
rect 287060 510614 287112 510620
rect 284300 484424 284352 484430
rect 284300 484366 284352 484372
rect 280068 461304 280120 461310
rect 280068 461246 280120 461252
rect 278688 461236 278740 461242
rect 278688 461178 278740 461184
rect 273996 461168 274048 461174
rect 273996 461110 274048 461116
rect 266360 460148 266412 460154
rect 266360 460090 266412 460096
rect 255044 458516 255096 458522
rect 255044 458458 255096 458464
rect 245568 458448 245620 458454
rect 245568 458390 245620 458396
rect 240784 458380 240836 458386
rect 240784 458322 240836 458328
rect 235908 458312 235960 458318
rect 235908 458254 235960 458260
rect 235920 457994 235948 458254
rect 240796 457994 240824 458322
rect 245580 457994 245608 458390
rect 255056 457994 255084 458458
rect 272016 458280 272072 458289
rect 272016 458215 272072 458224
rect 235796 457966 235948 457994
rect 240488 457966 240824 457994
rect 245272 457966 245608 457994
rect 254748 457966 255084 457994
rect 272030 457980 272058 458215
rect 274008 457994 274036 461110
rect 275560 458788 275612 458794
rect 275560 458730 275612 458736
rect 275572 457994 275600 458730
rect 277124 458720 277176 458726
rect 277124 458662 277176 458668
rect 277136 457994 277164 458662
rect 278700 457994 278728 461178
rect 280080 457994 280108 461246
rect 273700 457966 274036 457994
rect 275264 457966 275600 457994
rect 276828 457966 277164 457994
rect 278392 457966 278728 457994
rect 279956 457966 280108 457994
rect 284312 457994 284340 484366
rect 287072 480254 287100 510614
rect 288452 480254 288480 536794
rect 289820 524476 289872 524482
rect 289820 524418 289872 524424
rect 289832 480254 289860 524418
rect 287072 480226 287468 480254
rect 288452 480226 289032 480254
rect 289832 480226 290596 480254
rect 285864 470620 285916 470626
rect 285864 470562 285916 470568
rect 285876 457994 285904 470562
rect 287440 457994 287468 480226
rect 289004 457994 289032 480226
rect 290568 457994 290596 480226
rect 292592 457994 292620 563042
rect 293972 457994 294000 590650
rect 295340 576904 295392 576910
rect 295340 576846 295392 576852
rect 295352 457994 295380 576846
rect 296732 480254 296760 616830
rect 298112 480254 298140 643078
rect 296732 480226 296944 480254
rect 298112 480226 298508 480254
rect 296916 457994 296944 480226
rect 298480 457994 298508 480226
rect 299492 465730 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 328460 700800 328512 700806
rect 328460 700742 328512 700748
rect 318800 700732 318852 700738
rect 318800 700674 318852 700680
rect 303620 696992 303672 696998
rect 303620 696934 303672 696940
rect 300860 670812 300912 670818
rect 300860 670754 300912 670760
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299584 480254 299612 630634
rect 300872 480254 300900 670754
rect 299584 480226 300072 480254
rect 300872 480226 301728 480254
rect 299480 465724 299532 465730
rect 299480 465666 299532 465672
rect 300044 457994 300072 480226
rect 301700 457994 301728 480226
rect 303632 457994 303660 696934
rect 305000 683188 305052 683194
rect 305000 683130 305052 683136
rect 305012 457994 305040 683130
rect 306380 660340 306432 660346
rect 306380 660282 306432 660288
rect 306392 457994 306420 660282
rect 318812 480254 318840 700674
rect 320180 527876 320232 527882
rect 320180 527818 320232 527824
rect 320192 480254 320220 527818
rect 318812 480226 319024 480254
rect 320192 480226 320680 480254
rect 316040 464364 316092 464370
rect 316040 464306 316092 464312
rect 311808 461644 311860 461650
rect 311808 461586 311860 461592
rect 308680 460556 308732 460562
rect 308680 460498 308732 460504
rect 308692 457994 308720 460498
rect 310244 460488 310296 460494
rect 310244 460430 310296 460436
rect 310256 457994 310284 460430
rect 311820 457994 311848 461586
rect 313096 460760 313148 460766
rect 313096 460702 313148 460708
rect 284312 457966 284740 457994
rect 285876 457966 286304 457994
rect 287440 457966 287868 457994
rect 289004 457966 289432 457994
rect 290568 457966 290996 457994
rect 292592 457966 292652 457994
rect 293972 457966 294216 457994
rect 295352 457966 295780 457994
rect 296916 457966 297344 457994
rect 298480 457966 298908 457994
rect 300044 457966 300472 457994
rect 301700 457966 302128 457994
rect 303632 457966 303692 457994
rect 305012 457966 305256 457994
rect 306392 457966 306820 457994
rect 308384 457966 308720 457994
rect 309948 457966 310284 457994
rect 311604 457966 311848 457994
rect 313108 457858 313136 460702
rect 315028 460692 315080 460698
rect 315028 460634 315080 460640
rect 315040 457994 315068 460634
rect 314732 457966 315068 457994
rect 316052 457994 316080 464306
rect 318156 460896 318208 460902
rect 318156 460838 318208 460844
rect 318168 457994 318196 460838
rect 316052 457966 316296 457994
rect 317860 457966 318196 457994
rect 318996 457994 319024 480226
rect 320652 457994 320680 480226
rect 325700 465724 325752 465730
rect 325700 465666 325752 465672
rect 324136 460080 324188 460086
rect 324136 460022 324188 460028
rect 322848 460012 322900 460018
rect 322848 459954 322900 459960
rect 322860 457994 322888 459954
rect 318996 457966 319424 457994
rect 320652 457966 321080 457994
rect 322644 457966 322888 457994
rect 324148 457858 324176 460022
rect 325712 457994 325740 465666
rect 327080 460148 327132 460154
rect 327080 460090 327132 460096
rect 327092 457994 327120 460090
rect 328472 457994 328500 700742
rect 329840 698964 329892 698970
rect 329840 698906 329892 698912
rect 329852 480254 329880 698906
rect 329852 480226 330156 480254
rect 330128 457994 330156 480226
rect 331232 460018 331260 702986
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332600 700664 332652 700670
rect 332600 700606 332652 700612
rect 332612 480254 332640 700606
rect 338120 700596 338172 700602
rect 338120 700538 338172 700544
rect 332612 480226 333284 480254
rect 331772 460828 331824 460834
rect 331772 460770 331824 460776
rect 331220 460012 331272 460018
rect 331220 459954 331272 459960
rect 331784 457994 331812 460770
rect 333256 457994 333284 480226
rect 334808 467152 334860 467158
rect 334808 467094 334860 467100
rect 334820 457994 334848 467094
rect 336740 460624 336792 460630
rect 336740 460566 336792 460572
rect 336752 457994 336780 460566
rect 338132 457994 338160 700538
rect 342260 700528 342312 700534
rect 342260 700470 342312 700476
rect 340880 700460 340932 700466
rect 340880 700402 340932 700408
rect 340892 480254 340920 700402
rect 342272 480254 342300 700470
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 345032 480254 345060 700266
rect 340892 480226 341196 480254
rect 342272 480226 342760 480254
rect 345032 480226 345888 480254
rect 339592 468512 339644 468518
rect 339592 468454 339644 468460
rect 339604 457994 339632 468454
rect 341168 457994 341196 480226
rect 342732 457994 342760 480226
rect 344374 460320 344430 460329
rect 344374 460255 344430 460264
rect 344388 457994 344416 460255
rect 345860 457994 345888 480226
rect 347792 460086 347820 702406
rect 347872 700392 347924 700398
rect 347872 700334 347924 700340
rect 347780 460080 347832 460086
rect 347780 460022 347832 460028
rect 347884 458266 347912 700334
rect 351920 670744 351972 670750
rect 351920 670686 351972 670692
rect 350540 656940 350592 656946
rect 350540 656882 350592 656888
rect 350552 480254 350580 656882
rect 351932 480254 351960 670686
rect 356060 618316 356112 618322
rect 356060 618258 356112 618264
rect 354680 605872 354732 605878
rect 354680 605814 354732 605820
rect 354692 480254 354720 605814
rect 356072 480254 356100 618258
rect 361580 565888 361632 565894
rect 361580 565830 361632 565836
rect 360200 553444 360252 553450
rect 360200 553386 360252 553392
rect 350552 480226 350672 480254
rect 351932 480226 352236 480254
rect 354692 480226 355364 480254
rect 356072 480226 356928 480254
rect 349158 460184 349214 460193
rect 349158 460119 349214 460128
rect 347838 458238 347912 458266
rect 325712 457966 325772 457994
rect 327092 457966 327336 457994
rect 328472 457966 328900 457994
rect 330128 457966 330556 457994
rect 331784 457966 332120 457994
rect 333256 457966 333684 457994
rect 334820 457966 335248 457994
rect 336752 457966 336812 457994
rect 338132 457966 338376 457994
rect 339604 457966 340032 457994
rect 341168 457966 341596 457994
rect 342732 457966 343160 457994
rect 344388 457966 344724 457994
rect 345860 457966 346288 457994
rect 347838 457980 347866 458238
rect 349172 457994 349200 460119
rect 350644 457994 350672 480226
rect 352208 457994 352236 480226
rect 353852 460420 353904 460426
rect 353852 460362 353904 460368
rect 353864 457994 353892 460362
rect 355336 457994 355364 480226
rect 355968 459604 356020 459610
rect 355968 459546 356020 459552
rect 349172 457966 349508 457994
rect 350644 457966 351072 457994
rect 352208 457966 352636 457994
rect 353864 457966 354200 457994
rect 355336 457966 355764 457994
rect 313108 457830 313168 457858
rect 324148 457830 324208 457858
rect 281632 457632 281684 457638
rect 281520 457580 281632 457586
rect 281520 457574 281684 457580
rect 281520 457558 281672 457574
rect 355980 457502 356008 459546
rect 356900 457994 356928 480226
rect 358820 460352 358872 460358
rect 358820 460294 358872 460300
rect 358832 457994 358860 460294
rect 360212 457994 360240 553386
rect 361592 480254 361620 565830
rect 364352 527882 364380 702406
rect 364340 527876 364392 527882
rect 364340 527818 364392 527824
rect 365720 514820 365772 514826
rect 365720 514762 365772 514768
rect 364340 501016 364392 501022
rect 364340 500958 364392 500964
rect 364352 480254 364380 500958
rect 365732 480254 365760 514762
rect 361592 480226 361712 480254
rect 364352 480226 364840 480254
rect 365732 480226 366404 480254
rect 361684 457994 361712 480226
rect 363328 460284 363380 460290
rect 363328 460226 363380 460232
rect 363340 457994 363368 460226
rect 364812 457994 364840 480226
rect 366376 457994 366404 480226
rect 375932 462528 375984 462534
rect 375932 462470 375984 462476
rect 371240 462392 371292 462398
rect 371240 462334 371292 462340
rect 369860 461372 369912 461378
rect 369860 461314 369912 461320
rect 368112 460216 368164 460222
rect 368112 460158 368164 460164
rect 368124 457994 368152 460158
rect 369872 457994 369900 461314
rect 371252 457994 371280 462334
rect 374368 459604 374420 459610
rect 374368 459546 374420 459552
rect 373126 458244 373178 458250
rect 373126 458186 373178 458192
rect 356900 457966 357328 457994
rect 358832 457966 358984 457994
rect 360212 457966 360548 457994
rect 361684 457966 362112 457994
rect 363340 457966 363676 457994
rect 364812 457966 365240 457994
rect 366376 457966 366804 457994
rect 368124 457966 368460 457994
rect 369872 457966 370024 457994
rect 371252 457966 371588 457994
rect 373138 457980 373166 458186
rect 374380 457994 374408 459546
rect 375944 457994 375972 462470
rect 380900 462460 380952 462466
rect 380900 462402 380952 462408
rect 379152 461100 379204 461106
rect 379152 461042 379204 461048
rect 377588 458856 377640 458862
rect 377588 458798 377640 458804
rect 377600 457994 377628 458798
rect 379164 457994 379192 461042
rect 380912 457994 380940 462402
rect 396540 461032 396592 461038
rect 396540 460974 396592 460980
rect 391940 460964 391992 460970
rect 391940 460906 391992 460912
rect 382280 458652 382332 458658
rect 382280 458594 382332 458600
rect 382292 457994 382320 458594
rect 387064 458584 387116 458590
rect 387064 458526 387116 458532
rect 387076 457994 387104 458526
rect 391952 457994 391980 460906
rect 396552 457994 396580 460974
rect 397472 460902 397500 703520
rect 413664 700738 413692 703520
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 429212 464370 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 460204 700324 460256 700330
rect 460204 700266 460256 700272
rect 460216 660346 460244 700266
rect 460204 660340 460256 660346
rect 460204 660282 460256 660288
rect 429200 464364 429252 464370
rect 429200 464306 429252 464312
rect 417516 461304 417568 461310
rect 417516 461246 417568 461252
rect 397460 460896 397512 460902
rect 397460 460838 397512 460844
rect 407578 459776 407634 459785
rect 407578 459711 407634 459720
rect 407592 457994 407620 459711
rect 417424 458380 417476 458386
rect 417424 458322 417476 458328
rect 374380 457966 374716 457994
rect 375944 457966 376280 457994
rect 377600 457966 377936 457994
rect 379164 457966 379500 457994
rect 380912 457966 381064 457994
rect 382292 457966 382628 457994
rect 387076 457966 387412 457994
rect 391952 457966 392104 457994
rect 396552 457966 396888 457994
rect 407592 457966 407928 457994
rect 283380 457496 283432 457502
rect 237654 457464 237710 457473
rect 237360 457422 237654 457450
rect 239218 457464 239274 457473
rect 238924 457422 239218 457450
rect 237654 457399 237710 457408
rect 242346 457464 242402 457473
rect 242052 457422 242346 457450
rect 239218 457399 239274 457408
rect 243910 457464 243966 457473
rect 243616 457422 243910 457450
rect 242346 457399 242402 457408
rect 243910 457399 243966 457408
rect 246670 457464 246726 457473
rect 248234 457464 248290 457473
rect 246726 457422 246836 457450
rect 246670 457399 246726 457408
rect 250258 457464 250314 457473
rect 248290 457422 248400 457450
rect 249964 457422 250258 457450
rect 248234 457399 248290 457408
rect 251822 457464 251878 457473
rect 251528 457422 251822 457450
rect 250258 457399 250314 457408
rect 253386 457464 253442 457473
rect 253092 457422 253386 457450
rect 251822 457399 251878 457408
rect 256514 457464 256570 457473
rect 256312 457422 256514 457450
rect 253386 457399 253442 457408
rect 256514 457399 256570 457408
rect 257710 457464 257766 457473
rect 259274 457464 259330 457473
rect 257766 457422 257876 457450
rect 257710 457399 257766 457408
rect 261298 457464 261354 457473
rect 259330 457422 259440 457450
rect 261004 457422 261298 457450
rect 259274 457399 259330 457408
rect 262862 457464 262918 457473
rect 262568 457422 262862 457450
rect 261298 457399 261354 457408
rect 264518 457464 264574 457473
rect 264224 457422 264518 457450
rect 262862 457399 262918 457408
rect 266082 457464 266138 457473
rect 265788 457422 266082 457450
rect 264518 457399 264574 457408
rect 267554 457464 267610 457473
rect 267352 457422 267554 457450
rect 266082 457399 266138 457408
rect 267554 457399 267610 457408
rect 268750 457464 268806 457473
rect 270590 457464 270646 457473
rect 268806 457422 268916 457450
rect 270480 457422 270590 457450
rect 268750 457399 268806 457408
rect 283176 457444 283380 457450
rect 283176 457438 283432 457444
rect 355968 457496 356020 457502
rect 355968 457438 356020 457444
rect 383842 457464 383898 457473
rect 283176 457422 283420 457438
rect 270590 457399 270646 457408
rect 385406 457464 385462 457473
rect 383898 457422 384192 457450
rect 383842 457399 383898 457408
rect 388626 457464 388682 457473
rect 385462 457422 385756 457450
rect 385406 457399 385462 457408
rect 390190 457464 390246 457473
rect 388682 457422 388976 457450
rect 388626 457399 388682 457408
rect 393502 457464 393558 457473
rect 390246 457422 390540 457450
rect 390190 457399 390246 457408
rect 394882 457464 394938 457473
rect 393558 457422 393668 457450
rect 393502 457399 393558 457408
rect 398102 457464 398158 457473
rect 394938 457422 395232 457450
rect 394882 457399 394938 457408
rect 399666 457464 399722 457473
rect 398158 457422 398452 457450
rect 398102 457399 398158 457408
rect 401230 457464 401286 457473
rect 399722 457422 400016 457450
rect 399666 457399 399722 457408
rect 402978 457464 403034 457473
rect 401286 457422 401580 457450
rect 401230 457399 401286 457408
rect 404358 457464 404414 457473
rect 403034 457422 403144 457450
rect 402978 457399 403034 457408
rect 406014 457464 406070 457473
rect 404414 457422 404708 457450
rect 404358 457399 404414 457408
rect 409142 457464 409198 457473
rect 406070 457422 406364 457450
rect 406014 457399 406070 457408
rect 410706 457464 410762 457473
rect 409198 457422 409492 457450
rect 409142 457399 409198 457408
rect 412270 457464 412326 457473
rect 410762 457422 411056 457450
rect 410706 457399 410762 457408
rect 412326 457422 412620 457450
rect 414184 457422 414980 457450
rect 412270 457399 412326 457408
rect 233976 449880 234028 449886
rect 233976 449822 234028 449828
rect 233884 372564 233936 372570
rect 233884 372506 233936 372512
rect 309212 338150 309456 338178
rect 234816 338014 235152 338042
rect 235276 338014 235428 338042
rect 235552 338014 235796 338042
rect 236104 338014 236164 338042
rect 236288 338014 236532 338042
rect 236656 338014 236900 338042
rect 237024 338014 237268 338042
rect 237484 338014 237636 338042
rect 237760 338014 238004 338042
rect 238128 338014 238372 338042
rect 238496 338014 238740 338042
rect 238956 338014 239108 338042
rect 239232 338014 239476 338042
rect 239600 338014 239844 338042
rect 240152 338014 240212 338042
rect 240336 338014 240580 338042
rect 240704 338014 240948 338042
rect 241072 338014 241316 338042
rect 233976 336728 234028 336734
rect 233976 336670 234028 336676
rect 233884 336456 233936 336462
rect 233884 336398 233936 336404
rect 232504 320136 232556 320142
rect 232504 320078 232556 320084
rect 232594 319424 232650 319433
rect 232594 319359 232650 319368
rect 231860 275392 231912 275398
rect 231860 275334 231912 275340
rect 231124 267708 231176 267714
rect 231124 267650 231176 267656
rect 230480 240780 230532 240786
rect 230480 240722 230532 240728
rect 229744 164212 229796 164218
rect 229744 164154 229796 164160
rect 230492 16574 230520 240722
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227536 11688 227588 11694
rect 227536 11630 227588 11636
rect 226352 6886 226472 6914
rect 226352 480 226380 6886
rect 227548 480 227576 11630
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 275334
rect 232608 241466 232636 319359
rect 233240 247784 233292 247790
rect 233240 247726 233292 247732
rect 232596 241460 232648 241466
rect 232596 241402 232648 241408
rect 233252 16574 233280 247726
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 233896 4826 233924 336398
rect 233988 247722 234016 336670
rect 234620 330472 234672 330478
rect 234620 330414 234672 330420
rect 233976 247716 234028 247722
rect 233976 247658 234028 247664
rect 234632 49026 234660 330414
rect 234816 326398 234844 338014
rect 234804 326392 234856 326398
rect 234804 326334 234856 326340
rect 235276 316034 235304 338014
rect 235552 330478 235580 338014
rect 235540 330472 235592 330478
rect 235540 330414 235592 330420
rect 234724 316006 235304 316034
rect 234724 275330 234752 316006
rect 236104 283626 236132 338014
rect 236288 336054 236316 338014
rect 236276 336048 236328 336054
rect 236276 335990 236328 335996
rect 236656 316034 236684 338014
rect 237024 336734 237052 338014
rect 237012 336728 237064 336734
rect 237012 336670 237064 336676
rect 236196 316006 236684 316034
rect 236092 283620 236144 283626
rect 236092 283562 236144 283568
rect 234712 275324 234764 275330
rect 234712 275266 234764 275272
rect 234620 49020 234672 49026
rect 234620 48962 234672 48968
rect 234620 17400 234672 17406
rect 234620 17342 234672 17348
rect 233884 4820 233936 4826
rect 233884 4762 233936 4768
rect 234632 3194 234660 17342
rect 234712 6248 234764 6254
rect 234712 6190 234764 6196
rect 234620 3188 234672 3194
rect 234620 3130 234672 3136
rect 234724 1714 234752 6190
rect 236196 3369 236224 316006
rect 237484 11762 237512 338014
rect 237760 335354 237788 338014
rect 238128 336122 238156 338014
rect 238116 336116 238168 336122
rect 238116 336058 238168 336064
rect 237576 335326 237788 335354
rect 237576 203590 237604 335326
rect 238496 316034 238524 338014
rect 238760 330676 238812 330682
rect 238760 330618 238812 330624
rect 237668 316006 238524 316034
rect 237564 203584 237616 203590
rect 237564 203526 237616 203532
rect 237564 44872 237616 44878
rect 237564 44814 237616 44820
rect 237472 11756 237524 11762
rect 237472 11698 237524 11704
rect 237012 7676 237064 7682
rect 237012 7618 237064 7624
rect 236182 3360 236238 3369
rect 236182 3295 236238 3304
rect 235816 3188 235868 3194
rect 235816 3130 235868 3136
rect 234632 1686 234752 1714
rect 234632 480 234660 1686
rect 235828 480 235856 3130
rect 237024 480 237052 7618
rect 237576 6914 237604 44814
rect 237668 16574 237696 316006
rect 237668 16546 237788 16574
rect 237576 6886 237696 6914
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 354 237696 6886
rect 237760 6186 237788 16546
rect 237748 6180 237800 6186
rect 237748 6122 237800 6128
rect 238772 3505 238800 330618
rect 238852 330540 238904 330546
rect 238852 330482 238904 330488
rect 238864 18630 238892 330482
rect 238956 213246 238984 338014
rect 239232 330546 239260 338014
rect 239404 336728 239456 336734
rect 239404 336670 239456 336676
rect 239220 330540 239272 330546
rect 239220 330482 239272 330488
rect 239416 280838 239444 336670
rect 239600 330682 239628 338014
rect 240152 336734 240180 338014
rect 240140 336728 240192 336734
rect 240140 336670 240192 336676
rect 239588 330676 239640 330682
rect 239588 330618 239640 330624
rect 240232 330540 240284 330546
rect 240232 330482 240284 330488
rect 239404 280832 239456 280838
rect 239404 280774 239456 280780
rect 238944 213240 238996 213246
rect 238944 213182 238996 213188
rect 238852 18624 238904 18630
rect 238852 18566 238904 18572
rect 238944 18624 238996 18630
rect 238944 18566 238996 18572
rect 238956 16574 238984 18566
rect 238956 16546 239352 16574
rect 238758 3496 238814 3505
rect 238758 3431 238814 3440
rect 239324 480 239352 16546
rect 240244 3466 240272 330482
rect 240336 253230 240364 338014
rect 240704 330546 240732 338014
rect 240692 330540 240744 330546
rect 240692 330482 240744 330488
rect 241072 316034 241100 338014
rect 241670 337770 241698 338028
rect 241808 338014 242052 338042
rect 242176 338014 242420 338042
rect 242544 338014 242788 338042
rect 242912 338014 243156 338042
rect 243280 338014 243524 338042
rect 243648 338014 243892 338042
rect 244016 338014 244260 338042
rect 244384 338014 244628 338042
rect 244752 338014 244996 338042
rect 245120 338014 245364 338042
rect 245732 338014 245884 338042
rect 241670 337742 241744 337770
rect 241520 330540 241572 330546
rect 241520 330482 241572 330488
rect 240428 316006 241100 316034
rect 240324 253224 240376 253230
rect 240324 253166 240376 253172
rect 240324 26920 240376 26926
rect 240324 26862 240376 26868
rect 240232 3460 240284 3466
rect 240232 3402 240284 3408
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240336 354 240364 26862
rect 240428 3534 240456 316006
rect 241532 3602 241560 330482
rect 241612 329724 241664 329730
rect 241612 329666 241664 329672
rect 241624 3670 241652 329666
rect 241716 250510 241744 337742
rect 241808 302938 241836 338014
rect 242176 330546 242204 338014
rect 242164 330540 242216 330546
rect 242164 330482 242216 330488
rect 242544 329730 242572 338014
rect 242532 329724 242584 329730
rect 242532 329666 242584 329672
rect 242912 329118 242940 338014
rect 243280 335354 243308 338014
rect 243004 335326 243308 335354
rect 242900 329112 242952 329118
rect 242900 329054 242952 329060
rect 241796 302932 241848 302938
rect 241796 302874 241848 302880
rect 241704 250504 241756 250510
rect 241704 250446 241756 250452
rect 243004 206310 243032 335326
rect 243084 330540 243136 330546
rect 243084 330482 243136 330488
rect 243096 251870 243124 330482
rect 243648 316034 243676 338014
rect 244016 330546 244044 338014
rect 244004 330540 244056 330546
rect 244004 330482 244056 330488
rect 244280 326392 244332 326398
rect 244280 326334 244332 326340
rect 243188 316006 243676 316034
rect 243084 251864 243136 251870
rect 243084 251806 243136 251812
rect 242992 206304 243044 206310
rect 242992 206246 243044 206252
rect 241704 46232 241756 46238
rect 241704 46174 241756 46180
rect 241612 3664 241664 3670
rect 241612 3606 241664 3612
rect 241520 3596 241572 3602
rect 241520 3538 241572 3544
rect 240416 3528 240468 3534
rect 240416 3470 240468 3476
rect 241716 480 241744 46174
rect 242992 28280 243044 28286
rect 242992 28222 243044 28228
rect 243004 16574 243032 28222
rect 243004 16546 243124 16574
rect 242900 6180 242952 6186
rect 242900 6122 242952 6128
rect 242912 480 242940 6122
rect 243096 3482 243124 16546
rect 243188 3738 243216 316006
rect 244292 3806 244320 326334
rect 244384 204950 244412 338014
rect 244752 326398 244780 338014
rect 245120 336682 245148 338014
rect 244844 336654 245148 336682
rect 244740 326392 244792 326398
rect 244740 326334 244792 326340
rect 244844 316034 244872 336654
rect 244924 335572 244976 335578
rect 244924 335514 244976 335520
rect 244476 316006 244872 316034
rect 244476 221474 244504 316006
rect 244936 289134 244964 335514
rect 245752 326392 245804 326398
rect 245752 326334 245804 326340
rect 244924 289128 244976 289134
rect 244924 289070 244976 289076
rect 244464 221468 244516 221474
rect 244464 221410 244516 221416
rect 244372 204944 244424 204950
rect 244372 204886 244424 204892
rect 244372 47592 244424 47598
rect 244372 47534 244424 47540
rect 244384 16574 244412 47534
rect 245764 21418 245792 326334
rect 245856 254590 245884 338014
rect 245948 338014 246100 338042
rect 246224 338014 246468 338042
rect 246592 338014 246836 338042
rect 245844 254584 245896 254590
rect 245844 254526 245896 254532
rect 245752 21412 245804 21418
rect 245752 21354 245804 21360
rect 244384 16546 245240 16574
rect 244280 3800 244332 3806
rect 244280 3742 244332 3748
rect 243176 3732 243228 3738
rect 243176 3674 243228 3680
rect 243096 3454 244136 3482
rect 244108 480 244136 3454
rect 245212 480 245240 16546
rect 245948 3874 245976 338014
rect 246224 335578 246252 338014
rect 246212 335572 246264 335578
rect 246212 335514 246264 335520
rect 246592 326398 246620 338014
rect 247098 337770 247126 338028
rect 247328 338014 247480 338042
rect 247604 338014 247848 338042
rect 247972 338014 248216 338042
rect 248432 338014 248584 338042
rect 248708 338014 248952 338042
rect 249076 338014 249320 338042
rect 249444 338014 249688 338042
rect 249996 338014 250056 338042
rect 250180 338014 250424 338042
rect 250548 338014 250792 338042
rect 250916 338014 251160 338042
rect 251284 338014 251528 338042
rect 251652 338014 251896 338042
rect 252020 338014 252264 338042
rect 247098 337742 247172 337770
rect 246580 326392 246632 326398
rect 246580 326334 246632 326340
rect 247040 326392 247092 326398
rect 247040 326334 247092 326340
rect 246396 4820 246448 4826
rect 246396 4762 246448 4768
rect 245936 3868 245988 3874
rect 245936 3810 245988 3816
rect 246408 480 246436 4762
rect 247052 4010 247080 326334
rect 247040 4004 247092 4010
rect 247040 3946 247092 3952
rect 247144 3942 247172 337742
rect 247328 324970 247356 338014
rect 247604 335354 247632 338014
rect 247420 335326 247632 335354
rect 247316 324964 247368 324970
rect 247316 324906 247368 324912
rect 247420 321554 247448 335326
rect 247972 326398 248000 338014
rect 247960 326392 248012 326398
rect 247960 326334 248012 326340
rect 247236 321526 247448 321554
rect 247236 256018 247264 321526
rect 248432 320822 248460 338014
rect 248708 321554 248736 338014
rect 248524 321526 248736 321554
rect 248420 320816 248472 320822
rect 248420 320758 248472 320764
rect 247224 256012 247276 256018
rect 247224 255954 247276 255960
rect 248524 72486 248552 321526
rect 248604 320816 248656 320822
rect 248604 320758 248656 320764
rect 248616 220114 248644 320758
rect 249076 316034 249104 338014
rect 249444 331906 249472 338014
rect 249432 331900 249484 331906
rect 249432 331842 249484 331848
rect 249800 326392 249852 326398
rect 249800 326334 249852 326340
rect 248708 316006 249104 316034
rect 248604 220108 248656 220114
rect 248604 220050 248656 220056
rect 248512 72480 248564 72486
rect 248512 72422 248564 72428
rect 247224 29708 247276 29714
rect 247224 29650 247276 29656
rect 247236 16574 247264 29650
rect 248512 18692 248564 18698
rect 248512 18634 248564 18640
rect 247236 16546 247632 16574
rect 247132 3936 247184 3942
rect 247132 3878 247184 3884
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240336 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248524 354 248552 18634
rect 248708 4078 248736 316006
rect 249812 31074 249840 326334
rect 249892 326324 249944 326330
rect 249892 326266 249944 326272
rect 249904 217326 249932 326266
rect 249996 218754 250024 338014
rect 250180 326398 250208 338014
rect 250168 326392 250220 326398
rect 250168 326334 250220 326340
rect 250548 322250 250576 338014
rect 250916 326330 250944 338014
rect 251180 326392 251232 326398
rect 251180 326334 251232 326340
rect 250904 326324 250956 326330
rect 250904 326266 250956 326272
rect 250536 322244 250588 322250
rect 250536 322186 250588 322192
rect 249984 218748 250036 218754
rect 249984 218690 250036 218696
rect 249892 217320 249944 217326
rect 249892 217262 249944 217268
rect 251192 32434 251220 326334
rect 251284 64190 251312 338014
rect 251652 316034 251680 338014
rect 251824 335912 251876 335918
rect 251824 335854 251876 335860
rect 251376 316006 251680 316034
rect 251376 304298 251404 316006
rect 251364 304292 251416 304298
rect 251364 304234 251416 304240
rect 251836 215966 251864 335854
rect 252020 326398 252048 338014
rect 252618 337770 252646 338028
rect 252756 338014 253000 338042
rect 253124 338014 253368 338042
rect 253492 338014 253736 338042
rect 253952 338014 254104 338042
rect 254228 338014 254472 338042
rect 254596 338014 254840 338042
rect 254964 338014 255208 338042
rect 255516 338014 255576 338042
rect 255700 338014 255944 338042
rect 256068 338014 256312 338042
rect 256436 338014 256680 338042
rect 256896 338014 257048 338042
rect 257172 338014 257416 338042
rect 257540 338014 257784 338042
rect 258152 338014 258304 338042
rect 252618 337742 252692 337770
rect 252008 326392 252060 326398
rect 252008 326334 252060 326340
rect 251824 215960 251876 215966
rect 251824 215902 251876 215908
rect 252664 202162 252692 337742
rect 252756 330410 252784 338014
rect 253124 336818 253152 338014
rect 253032 336790 253152 336818
rect 253032 335918 253060 336790
rect 253492 336682 253520 338014
rect 253124 336654 253520 336682
rect 253020 335912 253072 335918
rect 253020 335854 253072 335860
rect 252744 330404 252796 330410
rect 252744 330346 252796 330352
rect 253124 316034 253152 336654
rect 253952 336598 253980 338014
rect 253204 336592 253256 336598
rect 253204 336534 253256 336540
rect 253940 336592 253992 336598
rect 253940 336534 253992 336540
rect 252756 316006 253152 316034
rect 252652 202156 252704 202162
rect 252652 202098 252704 202104
rect 251272 64184 251324 64190
rect 251272 64126 251324 64132
rect 251272 49020 251324 49026
rect 251272 48962 251324 48968
rect 251180 32428 251232 32434
rect 251180 32370 251232 32376
rect 249800 31068 249852 31074
rect 249800 31010 249852 31016
rect 251180 31068 251232 31074
rect 251180 31010 251232 31016
rect 249984 9172 250036 9178
rect 249984 9114 250036 9120
rect 248696 4072 248748 4078
rect 248696 4014 248748 4020
rect 249996 480 250024 9114
rect 251192 480 251220 31010
rect 251284 16574 251312 48962
rect 252756 29646 252784 316006
rect 253216 307086 253244 336534
rect 254228 335354 254256 338014
rect 254044 335326 254256 335354
rect 253204 307080 253256 307086
rect 253204 307022 253256 307028
rect 254044 284986 254072 335326
rect 254124 330540 254176 330546
rect 254124 330482 254176 330488
rect 254136 312594 254164 330482
rect 254596 316034 254624 338014
rect 254964 330546 254992 338014
rect 254952 330540 255004 330546
rect 254952 330482 255004 330488
rect 255412 330540 255464 330546
rect 255412 330482 255464 330488
rect 255320 330472 255372 330478
rect 255320 330414 255372 330420
rect 254228 316006 254624 316034
rect 254124 312588 254176 312594
rect 254124 312530 254176 312536
rect 254032 284980 254084 284986
rect 254032 284922 254084 284928
rect 254228 200802 254256 316006
rect 254216 200796 254268 200802
rect 254216 200738 254268 200744
rect 255332 61402 255360 330414
rect 255424 199442 255452 330482
rect 255516 214606 255544 338014
rect 255700 330546 255728 338014
rect 255688 330540 255740 330546
rect 255688 330482 255740 330488
rect 256068 316034 256096 338014
rect 256436 330478 256464 338014
rect 256700 330540 256752 330546
rect 256700 330482 256752 330488
rect 256424 330472 256476 330478
rect 256424 330414 256476 330420
rect 255608 316006 256096 316034
rect 255608 276690 255636 316006
rect 255596 276684 255648 276690
rect 255596 276626 255648 276632
rect 255504 214600 255556 214606
rect 255504 214542 255556 214548
rect 255412 199436 255464 199442
rect 255412 199378 255464 199384
rect 255320 61396 255372 61402
rect 255320 61338 255372 61344
rect 252744 29640 252796 29646
rect 252744 29582 252796 29588
rect 252560 21412 252612 21418
rect 252560 21354 252612 21360
rect 252572 16574 252600 21354
rect 255320 17332 255372 17338
rect 255320 17274 255372 17280
rect 255332 16574 255360 17274
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 254676 9104 254728 9110
rect 254676 9046 254728 9052
rect 254688 480 254716 9046
rect 255884 480 255912 16546
rect 256712 8974 256740 330482
rect 256792 330472 256844 330478
rect 256792 330414 256844 330420
rect 256804 33794 256832 330414
rect 256896 198014 256924 338014
rect 257172 330546 257200 338014
rect 257160 330540 257212 330546
rect 257160 330482 257212 330488
rect 257540 330478 257568 338014
rect 258276 330562 258304 338014
rect 258460 338014 258520 338042
rect 258644 338014 258888 338042
rect 259012 338014 259164 338042
rect 258172 330540 258224 330546
rect 258276 330534 258396 330562
rect 258172 330482 258224 330488
rect 257528 330472 257580 330478
rect 257528 330414 257580 330420
rect 258080 330336 258132 330342
rect 258080 330278 258132 330284
rect 256884 198008 256936 198014
rect 256884 197950 256936 197956
rect 256792 33788 256844 33794
rect 256792 33730 256844 33736
rect 256792 22840 256844 22846
rect 256792 22782 256844 22788
rect 256700 8968 256752 8974
rect 256700 8910 256752 8916
rect 248758 354 248870 480
rect 248524 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256804 354 256832 22782
rect 258092 9042 258120 330278
rect 258184 14482 258212 330482
rect 258264 330472 258316 330478
rect 258264 330414 258316 330420
rect 258276 196654 258304 330414
rect 258368 308446 258396 330534
rect 258460 330342 258488 338014
rect 258644 330546 258672 338014
rect 258632 330540 258684 330546
rect 258632 330482 258684 330488
rect 259012 330478 259040 338014
rect 259518 337770 259546 338028
rect 259656 338014 259900 338042
rect 260024 338014 260268 338042
rect 260392 338014 260636 338042
rect 259518 337742 259592 337770
rect 259460 330540 259512 330546
rect 259460 330482 259512 330488
rect 259000 330472 259052 330478
rect 259000 330414 259052 330420
rect 258448 330336 258500 330342
rect 258448 330278 258500 330284
rect 258356 308440 258408 308446
rect 258356 308382 258408 308388
rect 258264 196648 258316 196654
rect 258264 196590 258316 196596
rect 258264 32428 258316 32434
rect 258264 32370 258316 32376
rect 258172 14476 258224 14482
rect 258172 14418 258224 14424
rect 258080 9036 258132 9042
rect 258080 8978 258132 8984
rect 258276 480 258304 32370
rect 259472 10402 259500 330482
rect 259460 10396 259512 10402
rect 259460 10338 259512 10344
rect 259564 10334 259592 337742
rect 259656 14550 259684 338014
rect 260024 316034 260052 338014
rect 260392 330546 260420 338014
rect 260990 337770 261018 338028
rect 261128 338014 261372 338042
rect 261496 338014 261740 338042
rect 261864 338014 262108 338042
rect 262416 338014 262476 338042
rect 262600 338014 262844 338042
rect 262968 338014 263212 338042
rect 263336 338014 263580 338042
rect 263704 338014 263948 338042
rect 264072 338014 264316 338042
rect 264440 338014 264684 338042
rect 265052 338014 265204 338042
rect 260990 337742 261064 337770
rect 260840 336728 260892 336734
rect 260840 336670 260892 336676
rect 260380 330540 260432 330546
rect 260380 330482 260432 330488
rect 259748 316006 260052 316034
rect 259748 309806 259776 316006
rect 259736 309800 259788 309806
rect 259736 309742 259788 309748
rect 260852 55894 260880 336670
rect 260932 330540 260984 330546
rect 260932 330482 260984 330488
rect 260944 210458 260972 330482
rect 261036 211818 261064 337742
rect 261128 336734 261156 338014
rect 261116 336728 261168 336734
rect 261116 336670 261168 336676
rect 261496 316034 261524 338014
rect 261864 330546 261892 338014
rect 261852 330540 261904 330546
rect 261852 330482 261904 330488
rect 262220 330540 262272 330546
rect 262220 330482 262272 330488
rect 261128 316006 261524 316034
rect 261128 278050 261156 316006
rect 261116 278044 261168 278050
rect 261116 277986 261168 277992
rect 261024 211812 261076 211818
rect 261024 211754 261076 211760
rect 260932 210452 260984 210458
rect 260932 210394 260984 210400
rect 260840 55888 260892 55894
rect 260840 55830 260892 55836
rect 259736 19984 259788 19990
rect 259736 19926 259788 19932
rect 259644 14544 259696 14550
rect 259644 14486 259696 14492
rect 259552 10328 259604 10334
rect 259552 10270 259604 10276
rect 259748 6914 259776 19926
rect 260656 15972 260708 15978
rect 260656 15914 260708 15920
rect 259472 6886 259776 6914
rect 259472 480 259500 6886
rect 260668 480 260696 15914
rect 262232 14618 262260 330482
rect 262312 330472 262364 330478
rect 262312 330414 262364 330420
rect 262324 193866 262352 330414
rect 262416 195294 262444 338014
rect 262600 323610 262628 338014
rect 262968 330546 262996 338014
rect 262956 330540 263008 330546
rect 262956 330482 263008 330488
rect 263336 330478 263364 338014
rect 263704 336682 263732 338014
rect 263612 336654 263732 336682
rect 263324 330472 263376 330478
rect 263324 330414 263376 330420
rect 262588 323604 262640 323610
rect 262588 323546 262640 323552
rect 262404 195288 262456 195294
rect 262404 195230 262456 195236
rect 262312 193860 262364 193866
rect 262312 193802 262364 193808
rect 262312 25628 262364 25634
rect 262312 25570 262364 25576
rect 262324 16574 262352 25570
rect 262324 16546 262536 16574
rect 262220 14612 262272 14618
rect 262220 14554 262272 14560
rect 261760 10328 261812 10334
rect 261760 10270 261812 10276
rect 261772 480 261800 10270
rect 257038 354 257150 480
rect 256804 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 263612 13122 263640 336654
rect 264072 335354 264100 338014
rect 264440 336682 264468 338014
rect 263704 335326 264100 335354
rect 264164 336654 264468 336682
rect 263704 14686 263732 335326
rect 264164 316034 264192 336654
rect 264244 335980 264296 335986
rect 264244 335922 264296 335928
rect 263796 316006 264192 316034
rect 263796 192506 263824 316006
rect 264256 279478 264284 335922
rect 265072 330540 265124 330546
rect 265072 330482 265124 330488
rect 264244 279472 264296 279478
rect 264244 279414 264296 279420
rect 265084 222902 265112 330482
rect 265176 224262 265204 338014
rect 265268 338014 265420 338042
rect 265544 338014 265788 338042
rect 265912 338014 266156 338042
rect 265164 224256 265216 224262
rect 265164 224198 265216 224204
rect 265072 222896 265124 222902
rect 265072 222838 265124 222844
rect 263784 192500 263836 192506
rect 263784 192442 263836 192448
rect 263784 180124 263836 180130
rect 263784 180066 263836 180072
rect 263796 16574 263824 180066
rect 265268 60042 265296 338014
rect 265544 336190 265572 338014
rect 265532 336184 265584 336190
rect 265532 336126 265584 336132
rect 265912 330546 265940 338014
rect 266510 337770 266538 338028
rect 266648 338014 266892 338042
rect 267016 338014 267260 338042
rect 267384 338014 267628 338042
rect 267996 338014 268240 338042
rect 266510 337742 266584 337770
rect 265900 330540 265952 330546
rect 265900 330482 265952 330488
rect 266452 330540 266504 330546
rect 266452 330482 266504 330488
rect 266464 207670 266492 330482
rect 266556 209098 266584 337742
rect 266544 209092 266596 209098
rect 266544 209034 266596 209040
rect 266452 207664 266504 207670
rect 266452 207606 266504 207612
rect 265256 60036 265308 60042
rect 265256 59978 265308 59984
rect 264980 33788 265032 33794
rect 264980 33730 265032 33736
rect 263796 16546 264192 16574
rect 263692 14680 263744 14686
rect 263692 14622 263744 14628
rect 263600 13116 263652 13122
rect 263600 13058 263652 13064
rect 264164 480 264192 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 33730
rect 266648 4146 266676 338014
rect 267016 335986 267044 338014
rect 267004 335980 267056 335986
rect 267004 335922 267056 335928
rect 267384 330546 267412 338014
rect 267372 330540 267424 330546
rect 267372 330482 267424 330488
rect 267832 330540 267884 330546
rect 267832 330482 267884 330488
rect 267844 13190 267872 330482
rect 267924 329724 267976 329730
rect 267924 329666 267976 329672
rect 267936 14754 267964 329666
rect 268016 24200 268068 24206
rect 268016 24142 268068 24148
rect 267924 14748 267976 14754
rect 267924 14690 267976 14696
rect 267832 13184 267884 13190
rect 267832 13126 267884 13132
rect 266636 4140 266688 4146
rect 266636 4082 266688 4088
rect 268028 3602 268056 24142
rect 268108 14476 268160 14482
rect 268108 14418 268160 14424
rect 268016 3596 268068 3602
rect 268016 3538 268068 3544
rect 268120 3482 268148 14418
rect 266544 3460 266596 3466
rect 266544 3402 266596 3408
rect 267752 3454 268148 3482
rect 266556 480 266584 3402
rect 267752 480 267780 3454
rect 268212 3398 268240 338014
rect 268304 338014 268364 338042
rect 268488 338014 268732 338042
rect 268856 338014 269100 338042
rect 269224 338014 269468 338042
rect 269592 338014 269836 338042
rect 269960 338014 270204 338042
rect 268304 330546 268332 338014
rect 268292 330540 268344 330546
rect 268292 330482 268344 330488
rect 268488 329730 268516 338014
rect 268856 336258 268884 338014
rect 268844 336252 268896 336258
rect 268844 336194 268896 336200
rect 269120 330540 269172 330546
rect 269120 330482 269172 330488
rect 268476 329724 268528 329730
rect 268476 329666 268528 329672
rect 268476 3596 268528 3602
rect 268476 3538 268528 3544
rect 268200 3392 268252 3398
rect 268200 3334 268252 3340
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268488 354 268516 3538
rect 269132 3330 269160 330482
rect 269224 13258 269252 338014
rect 269304 336048 269356 336054
rect 269304 335990 269356 335996
rect 269316 329186 269344 335990
rect 269304 329180 269356 329186
rect 269304 329122 269356 329128
rect 269592 316034 269620 338014
rect 269764 336524 269816 336530
rect 269764 336466 269816 336472
rect 269316 316006 269620 316034
rect 269316 14822 269344 316006
rect 269776 286346 269804 336466
rect 269960 330546 269988 338014
rect 270558 337770 270586 338028
rect 270696 338014 270940 338042
rect 271064 338014 271216 338042
rect 271340 338014 271584 338042
rect 271892 338014 271952 338042
rect 272076 338014 272320 338042
rect 272444 338014 272688 338042
rect 272812 338014 273056 338042
rect 273272 338014 273424 338042
rect 273548 338014 273792 338042
rect 273916 338014 274160 338042
rect 274284 338014 274528 338042
rect 274836 338014 274896 338042
rect 275020 338014 275264 338042
rect 275388 338014 275632 338042
rect 275756 338014 276000 338042
rect 276124 338014 276368 338042
rect 276492 338014 276736 338042
rect 276860 338014 277104 338042
rect 277472 338014 277624 338042
rect 270558 337742 270632 337770
rect 269948 330540 270000 330546
rect 269948 330482 270000 330488
rect 269764 286340 269816 286346
rect 269764 286282 269816 286288
rect 269304 14816 269356 14822
rect 269304 14758 269356 14764
rect 270604 13326 270632 337742
rect 270696 15910 270724 338014
rect 271064 336326 271092 338014
rect 271144 336728 271196 336734
rect 271144 336670 271196 336676
rect 271052 336320 271104 336326
rect 271052 336262 271104 336268
rect 270776 330540 270828 330546
rect 270776 330482 270828 330488
rect 270684 15904 270736 15910
rect 270684 15846 270736 15852
rect 270788 13394 270816 330482
rect 271156 282198 271184 336670
rect 271340 330546 271368 338014
rect 271892 336530 271920 338014
rect 271880 336524 271932 336530
rect 271880 336466 271932 336472
rect 271328 330540 271380 330546
rect 271328 330482 271380 330488
rect 271972 330540 272024 330546
rect 271972 330482 272024 330488
rect 271984 316742 272012 330482
rect 271972 316736 272024 316742
rect 271972 316678 272024 316684
rect 271144 282192 271196 282198
rect 271144 282134 271196 282140
rect 270776 13388 270828 13394
rect 270776 13330 270828 13336
rect 270592 13320 270644 13326
rect 270592 13262 270644 13268
rect 269212 13252 269264 13258
rect 269212 13194 269264 13200
rect 270776 13116 270828 13122
rect 270776 13058 270828 13064
rect 270040 3528 270092 3534
rect 270040 3470 270092 3476
rect 269120 3324 269172 3330
rect 269120 3266 269172 3272
rect 270052 480 270080 3470
rect 268814 354 268926 480
rect 268488 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 13058
rect 271972 11756 272024 11762
rect 271972 11698 272024 11704
rect 271880 3596 271932 3602
rect 271880 3538 271932 3544
rect 271892 3262 271920 3538
rect 271984 3482 272012 11698
rect 272076 3602 272104 338014
rect 272444 336734 272472 338014
rect 272432 336728 272484 336734
rect 272432 336670 272484 336676
rect 272812 330546 272840 338014
rect 273272 336394 273300 338014
rect 273260 336388 273312 336394
rect 273260 336330 273312 336336
rect 273548 335354 273576 338014
rect 273916 336682 273944 338014
rect 273456 335326 273576 335354
rect 273824 336654 273944 336682
rect 272800 330540 272852 330546
rect 272800 330482 272852 330488
rect 273456 327758 273484 335326
rect 273444 327752 273496 327758
rect 273444 327694 273496 327700
rect 273352 326392 273404 326398
rect 273352 326334 273404 326340
rect 273364 35222 273392 326334
rect 273824 316034 273852 336654
rect 273904 335776 273956 335782
rect 273904 335718 273956 335724
rect 273548 316006 273852 316034
rect 273352 35216 273404 35222
rect 273352 35158 273404 35164
rect 273548 24138 273576 316006
rect 273916 287706 273944 335718
rect 274284 326398 274312 338014
rect 274272 326392 274324 326398
rect 274272 326334 274324 326340
rect 274640 326392 274692 326398
rect 274640 326334 274692 326340
rect 273904 287700 273956 287706
rect 273904 287642 273956 287648
rect 274652 273970 274680 326334
rect 274836 323678 274864 338014
rect 275020 326398 275048 338014
rect 275388 331214 275416 338014
rect 275112 331186 275416 331214
rect 275008 326392 275060 326398
rect 275008 326334 275060 326340
rect 274824 323672 274876 323678
rect 274824 323614 274876 323620
rect 275112 323490 275140 331186
rect 274744 323462 275140 323490
rect 274640 273964 274692 273970
rect 274640 273906 274692 273912
rect 274744 232558 274772 323462
rect 275756 321554 275784 338014
rect 276020 326392 276072 326398
rect 276020 326334 276072 326340
rect 274836 321526 275784 321554
rect 274836 308514 274864 321526
rect 274824 308508 274876 308514
rect 274824 308450 274876 308456
rect 274824 274100 274876 274106
rect 274824 274042 274876 274048
rect 274732 232552 274784 232558
rect 274732 232494 274784 232500
rect 273536 24132 273588 24138
rect 273536 24074 273588 24080
rect 272064 3596 272116 3602
rect 272064 3538 272116 3544
rect 273628 3596 273680 3602
rect 273628 3538 273680 3544
rect 271984 3454 272472 3482
rect 271880 3256 271932 3262
rect 271880 3198 271932 3204
rect 272444 480 272472 3454
rect 273640 480 273668 3538
rect 274836 480 274864 274042
rect 276032 43450 276060 326334
rect 276124 249082 276152 338014
rect 276492 326398 276520 338014
rect 276860 336682 276888 338014
rect 276584 336654 276888 336682
rect 276480 326392 276532 326398
rect 276480 326334 276532 326340
rect 276584 316034 276612 336654
rect 276664 336116 276716 336122
rect 276664 336058 276716 336064
rect 276676 325038 276704 336058
rect 277492 326392 277544 326398
rect 277492 326334 277544 326340
rect 276664 325032 276716 325038
rect 276664 324974 276716 324980
rect 276216 316006 276612 316034
rect 276216 309874 276244 316006
rect 276204 309868 276256 309874
rect 276204 309810 276256 309816
rect 276204 249212 276256 249218
rect 276204 249154 276256 249160
rect 276112 249076 276164 249082
rect 276112 249018 276164 249024
rect 276020 43444 276072 43450
rect 276020 43386 276072 43392
rect 276216 6914 276244 249154
rect 277504 246362 277532 326334
rect 277596 290494 277624 338014
rect 277688 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278576 338042
rect 278884 338014 278944 338042
rect 279068 338014 279312 338042
rect 279436 338014 279680 338042
rect 279804 338014 280048 338042
rect 277584 290488 277636 290494
rect 277584 290430 277636 290436
rect 277492 246356 277544 246362
rect 277492 246298 277544 246304
rect 277688 51746 277716 338014
rect 277964 335782 277992 338014
rect 277952 335776 278004 335782
rect 277952 335718 278004 335724
rect 278332 326398 278360 338014
rect 278320 326392 278372 326398
rect 278320 326334 278372 326340
rect 278780 326324 278832 326330
rect 278780 326266 278832 326272
rect 277676 51740 277728 51746
rect 277676 51682 277728 51688
rect 278792 22778 278820 326266
rect 278884 225622 278912 338014
rect 278964 326392 279016 326398
rect 278964 326334 279016 326340
rect 278976 244934 279004 326334
rect 279068 300150 279096 338014
rect 279436 326398 279464 338014
rect 279424 326392 279476 326398
rect 279424 326334 279476 326340
rect 279804 326330 279832 338014
rect 280402 337770 280430 338028
rect 280540 338014 280784 338042
rect 280908 338014 281152 338042
rect 281276 338014 281520 338042
rect 281644 338014 281888 338042
rect 282012 338014 282256 338042
rect 282380 338014 282624 338042
rect 282992 338014 283144 338042
rect 280402 337742 280476 337770
rect 280448 326534 280476 337742
rect 280436 326528 280488 326534
rect 280436 326470 280488 326476
rect 280252 326392 280304 326398
rect 280252 326334 280304 326340
rect 279792 326324 279844 326330
rect 279792 326266 279844 326272
rect 280160 323604 280212 323610
rect 280160 323546 280212 323552
rect 279056 300144 279108 300150
rect 279056 300086 279108 300092
rect 278964 244928 279016 244934
rect 278964 244870 279016 244876
rect 278872 225616 278924 225622
rect 278872 225558 278924 225564
rect 280172 50386 280200 323546
rect 280264 272542 280292 326334
rect 280540 321858 280568 338014
rect 280620 326528 280672 326534
rect 280620 326470 280672 326476
rect 280356 321830 280568 321858
rect 280356 291854 280384 321830
rect 280632 318794 280660 326470
rect 280908 323610 280936 338014
rect 281276 326398 281304 338014
rect 281264 326392 281316 326398
rect 281264 326334 281316 326340
rect 281540 326392 281592 326398
rect 281540 326334 281592 326340
rect 280896 323604 280948 323610
rect 280896 323546 280948 323552
rect 280448 318766 280660 318794
rect 280448 301510 280476 318766
rect 280436 301504 280488 301510
rect 280436 301446 280488 301452
rect 280344 291848 280396 291854
rect 280344 291790 280396 291796
rect 280252 272536 280304 272542
rect 280252 272478 280304 272484
rect 281552 53106 281580 326334
rect 281644 243574 281672 338014
rect 282012 326398 282040 338014
rect 282000 326392 282052 326398
rect 282000 326334 282052 326340
rect 282380 316034 282408 338014
rect 282920 328296 282972 328302
rect 282920 328238 282972 328244
rect 281736 316006 282408 316034
rect 281736 271182 281764 316006
rect 281724 271176 281776 271182
rect 281724 271118 281776 271124
rect 281632 243568 281684 243574
rect 281632 243510 281684 243516
rect 282932 71058 282960 328238
rect 283012 326936 283064 326942
rect 283012 326878 283064 326884
rect 283024 239426 283052 326878
rect 283116 242214 283144 338014
rect 283208 338014 283268 338042
rect 283392 338014 283636 338042
rect 283760 338014 284004 338042
rect 283208 328302 283236 338014
rect 283196 328296 283248 328302
rect 283196 328238 283248 328244
rect 283392 316034 283420 338014
rect 283760 326942 283788 338014
rect 284358 337770 284386 338028
rect 284496 338014 284740 338042
rect 284864 338014 285108 338042
rect 285232 338014 285476 338042
rect 285692 338014 285844 338042
rect 285968 338014 286212 338042
rect 286336 338014 286580 338042
rect 286704 338014 286948 338042
rect 287256 338014 287316 338042
rect 287440 338014 287684 338042
rect 287808 338014 288052 338042
rect 288176 338014 288420 338042
rect 288544 338014 288788 338042
rect 288912 338014 289156 338042
rect 289280 338014 289524 338042
rect 284358 337742 284432 337770
rect 283748 326936 283800 326942
rect 283748 326878 283800 326884
rect 283208 316006 283420 316034
rect 283208 303006 283236 316006
rect 283196 303000 283248 303006
rect 283196 302942 283248 302948
rect 283104 242208 283156 242214
rect 283104 242150 283156 242156
rect 283012 239420 283064 239426
rect 283012 239362 283064 239368
rect 282920 71052 282972 71058
rect 282920 70994 282972 71000
rect 284404 54534 284432 337742
rect 284496 336054 284524 338014
rect 284484 336048 284536 336054
rect 284484 335990 284536 335996
rect 284864 335354 284892 338014
rect 284496 335326 284892 335354
rect 284496 269822 284524 335326
rect 285232 316034 285260 338014
rect 285692 336122 285720 338014
rect 285680 336116 285732 336122
rect 285680 336058 285732 336064
rect 285772 330540 285824 330546
rect 285772 330482 285824 330488
rect 284588 316006 285260 316034
rect 284484 269816 284536 269822
rect 284484 269758 284536 269764
rect 284392 54528 284444 54534
rect 284392 54470 284444 54476
rect 281540 53100 281592 53106
rect 281540 53042 281592 53048
rect 280160 50380 280212 50386
rect 280160 50322 280212 50328
rect 284588 36582 284616 316006
rect 285680 284980 285732 284986
rect 285680 284922 285732 284928
rect 284576 36576 284628 36582
rect 284576 36518 284628 36524
rect 282920 35216 282972 35222
rect 282920 35158 282972 35164
rect 278780 22772 278832 22778
rect 278780 22714 278832 22720
rect 282932 16574 282960 35158
rect 285692 16574 285720 284922
rect 285784 238066 285812 330482
rect 285968 316034 285996 338014
rect 286232 336048 286284 336054
rect 286232 335990 286284 335996
rect 286244 325694 286272 335990
rect 286336 330546 286364 338014
rect 286416 336320 286468 336326
rect 286416 336262 286468 336268
rect 286324 330540 286376 330546
rect 286324 330482 286376 330488
rect 286244 325666 286364 325694
rect 285876 316006 285996 316034
rect 285876 268394 285904 316006
rect 286336 285054 286364 325666
rect 286428 312662 286456 336262
rect 286704 330614 286732 338014
rect 286692 330608 286744 330614
rect 286692 330550 286744 330556
rect 287152 330132 287204 330138
rect 287152 330074 287204 330080
rect 286416 312656 286468 312662
rect 286416 312598 286468 312604
rect 286324 285048 286376 285054
rect 286324 284990 286376 284996
rect 285864 268388 285916 268394
rect 285864 268330 285916 268336
rect 287164 264246 287192 330074
rect 287256 265674 287284 338014
rect 287440 316034 287468 338014
rect 287808 336326 287836 338014
rect 287796 336320 287848 336326
rect 287796 336262 287848 336268
rect 287704 335708 287756 335714
rect 287704 335650 287756 335656
rect 287348 316006 287468 316034
rect 287244 265668 287296 265674
rect 287244 265610 287296 265616
rect 287152 264240 287204 264246
rect 287152 264182 287204 264188
rect 285772 238060 285824 238066
rect 285772 238002 285824 238008
rect 287348 37942 287376 316006
rect 287716 289202 287744 335650
rect 288176 330138 288204 338014
rect 288164 330132 288216 330138
rect 288164 330074 288216 330080
rect 287704 289196 287756 289202
rect 287704 289138 287756 289144
rect 287336 37936 287388 37942
rect 287336 37878 287388 37884
rect 282932 16546 283144 16574
rect 285692 16546 286640 16574
rect 279056 15904 279108 15910
rect 279056 15846 279108 15852
rect 276032 6886 276244 6914
rect 276032 480 276060 6886
rect 278320 4888 278372 4894
rect 278320 4830 278372 4836
rect 277122 3360 277178 3369
rect 277122 3295 277178 3304
rect 277136 480 277164 3295
rect 278332 480 278360 4830
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 15846
rect 281908 6316 281960 6322
rect 281908 6258 281960 6264
rect 280712 3664 280764 3670
rect 280712 3606 280764 3612
rect 280724 480 280752 3606
rect 281920 480 281948 6258
rect 283116 480 283144 16546
rect 285404 4956 285456 4962
rect 285404 4898 285456 4904
rect 284300 3732 284352 3738
rect 284300 3674 284352 3680
rect 284312 480 284340 3674
rect 285416 480 285444 4898
rect 286612 480 286640 16546
rect 288544 10470 288572 338014
rect 288912 331974 288940 338014
rect 289280 336682 289308 338014
rect 289878 337770 289906 338028
rect 290016 338014 290260 338042
rect 290384 338014 290628 338042
rect 290752 338014 290996 338042
rect 291212 338014 291364 338042
rect 291488 338014 291732 338042
rect 291856 338014 292100 338042
rect 292224 338014 292468 338042
rect 292592 338014 292836 338042
rect 292960 338014 293204 338042
rect 293328 338014 293572 338042
rect 293696 338014 293940 338042
rect 294064 338014 294308 338042
rect 294432 338014 294676 338042
rect 294800 338014 295044 338042
rect 295168 338014 295320 338042
rect 295536 338014 295688 338042
rect 295812 338014 296056 338042
rect 296180 338014 296424 338042
rect 296732 338014 296792 338042
rect 296916 338014 297160 338042
rect 297284 338014 297528 338042
rect 297652 338014 297896 338042
rect 298204 338014 298264 338042
rect 298388 338014 298632 338042
rect 298756 338014 299000 338042
rect 299124 338014 299368 338042
rect 299676 338014 299736 338042
rect 299860 338014 300104 338042
rect 300228 338014 300472 338042
rect 300596 338014 300840 338042
rect 300964 338014 301208 338042
rect 301332 338014 301576 338042
rect 301700 338014 301944 338042
rect 302252 338014 302312 338042
rect 302436 338014 302680 338042
rect 302804 338014 303048 338042
rect 303172 338014 303416 338042
rect 303724 338014 303784 338042
rect 303908 338014 304152 338042
rect 304276 338014 304520 338042
rect 304644 338014 304888 338042
rect 305196 338014 305256 338042
rect 305380 338014 305624 338042
rect 305748 338014 305992 338042
rect 306116 338014 306360 338042
rect 306484 338014 306728 338042
rect 306852 338014 307096 338042
rect 307220 338014 307372 338042
rect 307496 338014 307740 338042
rect 307864 338014 308108 338042
rect 308232 338014 308476 338042
rect 308600 338014 308844 338042
rect 289878 337742 289952 337770
rect 289004 336654 289308 336682
rect 288900 331968 288952 331974
rect 288900 331910 288952 331916
rect 289004 316034 289032 336654
rect 289176 336592 289228 336598
rect 289176 336534 289228 336540
rect 289084 336116 289136 336122
rect 289084 336058 289136 336064
rect 288636 316006 289032 316034
rect 288532 10464 288584 10470
rect 288532 10406 288584 10412
rect 288636 7614 288664 316006
rect 288624 7608 288676 7614
rect 288624 7550 288676 7556
rect 288992 5024 289044 5030
rect 288992 4966 289044 4972
rect 287796 3800 287848 3806
rect 287796 3742 287848 3748
rect 287808 480 287836 3742
rect 289004 480 289032 4966
rect 289096 4826 289124 336058
rect 289188 286414 289216 336534
rect 289924 320890 289952 337742
rect 290016 336598 290044 338014
rect 290004 336592 290056 336598
rect 290004 336534 290056 336540
rect 290384 335714 290412 338014
rect 290372 335708 290424 335714
rect 290372 335650 290424 335656
rect 289912 320884 289964 320890
rect 289912 320826 289964 320832
rect 290752 316034 290780 338014
rect 291212 336054 291240 338014
rect 291200 336048 291252 336054
rect 291200 335990 291252 335996
rect 291488 335354 291516 338014
rect 291856 336682 291884 338014
rect 290016 316006 290780 316034
rect 291304 335326 291516 335354
rect 291672 336654 291884 336682
rect 289176 286408 289228 286414
rect 289176 286350 289228 286356
rect 290016 236706 290044 316006
rect 291304 262886 291332 335326
rect 291384 330540 291436 330546
rect 291384 330482 291436 330488
rect 291396 283694 291424 330482
rect 291672 316034 291700 336654
rect 291844 335980 291896 335986
rect 291844 335922 291896 335928
rect 291488 316006 291700 316034
rect 291384 283688 291436 283694
rect 291384 283630 291436 283636
rect 291292 262880 291344 262886
rect 291292 262822 291344 262828
rect 290004 236700 290056 236706
rect 290004 236642 290056 236648
rect 291488 40730 291516 316006
rect 291476 40724 291528 40730
rect 291476 40666 291528 40672
rect 291856 15978 291884 335922
rect 291936 335844 291988 335850
rect 291936 335786 291988 335792
rect 291948 322318 291976 335786
rect 292224 330546 292252 338014
rect 292212 330540 292264 330546
rect 292212 330482 292264 330488
rect 291936 322312 291988 322318
rect 291936 322254 291988 322260
rect 292592 320890 292620 338014
rect 292960 335354 292988 338014
rect 293224 336728 293276 336734
rect 293224 336670 293276 336676
rect 292868 335326 292988 335354
rect 292868 321554 292896 335326
rect 293236 326466 293264 336670
rect 293328 335850 293356 338014
rect 293316 335844 293368 335850
rect 293316 335786 293368 335792
rect 293224 326460 293276 326466
rect 293224 326402 293276 326408
rect 292684 321526 292896 321554
rect 292580 320884 292632 320890
rect 292580 320826 292632 320832
rect 292580 261588 292632 261594
rect 292580 261530 292632 261536
rect 292592 16574 292620 261530
rect 292684 235278 292712 321526
rect 292764 320884 292816 320890
rect 292764 320826 292816 320832
rect 292776 261526 292804 320826
rect 293696 316034 293724 338014
rect 292868 316006 293724 316034
rect 292764 261520 292816 261526
rect 292764 261462 292816 261468
rect 292868 260166 292896 316006
rect 292856 260160 292908 260166
rect 292856 260102 292908 260108
rect 292672 235272 292724 235278
rect 292672 235214 292724 235220
rect 294064 233918 294092 338014
rect 294432 336802 294460 338014
rect 294420 336796 294472 336802
rect 294420 336738 294472 336744
rect 294800 336682 294828 338014
rect 294156 336654 294828 336682
rect 294156 258738 294184 336654
rect 294604 336524 294656 336530
rect 294604 336466 294656 336472
rect 294236 326392 294288 326398
rect 294236 326334 294288 326340
rect 294144 258732 294196 258738
rect 294144 258674 294196 258680
rect 294052 233912 294104 233918
rect 294052 233854 294104 233860
rect 294248 42090 294276 326334
rect 294616 307154 294644 336466
rect 295168 326398 295196 338014
rect 295536 326466 295564 338014
rect 295812 335354 295840 338014
rect 295628 335326 295840 335354
rect 295984 335368 296036 335374
rect 295524 326460 295576 326466
rect 295524 326402 295576 326408
rect 295156 326392 295208 326398
rect 295156 326334 295208 326340
rect 295524 326256 295576 326262
rect 295524 326198 295576 326204
rect 295432 323604 295484 323610
rect 295432 323546 295484 323552
rect 295340 322108 295392 322114
rect 295340 322050 295392 322056
rect 294604 307148 294656 307154
rect 294604 307090 294656 307096
rect 294236 42084 294288 42090
rect 294236 42026 294288 42032
rect 295352 39370 295380 322050
rect 295444 257378 295472 323546
rect 295536 282266 295564 326198
rect 295628 323610 295656 335326
rect 295984 335310 296036 335316
rect 295616 323604 295668 323610
rect 295616 323546 295668 323552
rect 295524 282260 295576 282266
rect 295524 282202 295576 282208
rect 295996 280906 296024 335310
rect 296180 322114 296208 338014
rect 296732 335374 296760 338014
rect 296812 336728 296864 336734
rect 296812 336670 296864 336676
rect 296720 335368 296772 335374
rect 296720 335310 296772 335316
rect 296168 322108 296220 322114
rect 296168 322050 296220 322056
rect 295984 280900 296036 280906
rect 295984 280842 296036 280848
rect 296720 279676 296772 279682
rect 296720 279618 296772 279624
rect 295432 257372 295484 257378
rect 295432 257314 295484 257320
rect 295340 39364 295392 39370
rect 295340 39306 295392 39312
rect 296732 16574 296760 279618
rect 296824 231130 296852 336670
rect 296916 329254 296944 338014
rect 297284 336734 297312 338014
rect 297272 336728 297324 336734
rect 297272 336670 297324 336676
rect 297456 336456 297508 336462
rect 297456 336398 297508 336404
rect 297364 336184 297416 336190
rect 297364 336126 297416 336132
rect 296904 329248 296956 329254
rect 296904 329190 296956 329196
rect 296996 326392 297048 326398
rect 296996 326334 297048 326340
rect 297008 279546 297036 326334
rect 296996 279540 297048 279546
rect 296996 279482 297048 279488
rect 296812 231124 296864 231130
rect 296812 231066 296864 231072
rect 292592 16546 293264 16574
rect 296732 16546 297312 16574
rect 291844 15972 291896 15978
rect 291844 15914 291896 15920
rect 290188 7608 290240 7614
rect 290188 7550 290240 7556
rect 289084 4820 289136 4826
rect 289084 4762 289136 4768
rect 290200 480 290228 7550
rect 292580 4820 292632 4826
rect 292580 4762 292632 4768
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 291396 480 291424 3810
rect 292592 480 292620 4762
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 296076 5092 296128 5098
rect 296076 5034 296128 5040
rect 294880 3936 294932 3942
rect 294880 3878 294932 3884
rect 294892 480 294920 3878
rect 296088 480 296116 5034
rect 297284 480 297312 16546
rect 297376 9178 297404 336126
rect 297468 304366 297496 336398
rect 297652 326398 297680 338014
rect 297640 326392 297692 326398
rect 297640 326334 297692 326340
rect 297456 304360 297508 304366
rect 297456 304302 297508 304308
rect 298204 256086 298232 338014
rect 298388 335354 298416 338014
rect 298756 336818 298784 338014
rect 298572 336790 298784 336818
rect 298572 336530 298600 336790
rect 299124 336682 299152 338014
rect 298664 336654 299152 336682
rect 298560 336524 298612 336530
rect 298560 336466 298612 336472
rect 298296 335326 298416 335354
rect 298296 325106 298324 335326
rect 298284 325100 298336 325106
rect 298284 325042 298336 325048
rect 298664 316034 298692 336654
rect 298744 336592 298796 336598
rect 298744 336534 298796 336540
rect 298388 316006 298692 316034
rect 298192 256080 298244 256086
rect 298192 256022 298244 256028
rect 298388 254658 298416 316006
rect 298376 254652 298428 254658
rect 298376 254594 298428 254600
rect 298756 25566 298784 336534
rect 299572 326392 299624 326398
rect 299572 326334 299624 326340
rect 299480 253428 299532 253434
rect 299480 253370 299532 253376
rect 298744 25560 298796 25566
rect 298744 25502 298796 25508
rect 297364 9172 297416 9178
rect 297364 9114 297416 9120
rect 298468 4004 298520 4010
rect 298468 3946 298520 3952
rect 298480 480 298508 3946
rect 299492 2106 299520 253370
rect 299584 228410 299612 326334
rect 299676 229770 299704 338014
rect 299860 336462 299888 338014
rect 299848 336456 299900 336462
rect 299848 336398 299900 336404
rect 300228 316034 300256 338014
rect 300596 326398 300624 338014
rect 300768 336728 300820 336734
rect 300768 336670 300820 336676
rect 300780 334626 300808 336670
rect 300768 334620 300820 334626
rect 300768 334562 300820 334568
rect 300584 326392 300636 326398
rect 300584 326334 300636 326340
rect 300860 326392 300912 326398
rect 300860 326334 300912 326340
rect 299768 316006 300256 316034
rect 299768 253298 299796 316006
rect 299756 253292 299808 253298
rect 299756 253234 299808 253240
rect 299664 229764 299716 229770
rect 299664 229706 299716 229712
rect 299572 228404 299624 228410
rect 299572 228346 299624 228352
rect 300872 11830 300900 326334
rect 300964 278118 300992 338014
rect 301332 327826 301360 338014
rect 301504 335504 301556 335510
rect 301504 335446 301556 335452
rect 301320 327820 301372 327826
rect 301320 327762 301372 327768
rect 300952 278112 301004 278118
rect 300952 278054 301004 278060
rect 301516 18630 301544 335446
rect 301700 326398 301728 338014
rect 302252 336394 302280 338014
rect 302436 336598 302464 338014
rect 302424 336592 302476 336598
rect 302424 336534 302476 336540
rect 302240 336388 302292 336394
rect 302240 336330 302292 336336
rect 302332 330540 302384 330546
rect 302332 330482 302384 330488
rect 301688 326392 301740 326398
rect 301688 326334 301740 326340
rect 302344 276758 302372 330482
rect 302804 316034 302832 338014
rect 303068 336524 303120 336530
rect 303068 336466 303120 336472
rect 302884 336456 302936 336462
rect 302884 336398 302936 336404
rect 302436 316006 302832 316034
rect 302332 276752 302384 276758
rect 302332 276694 302384 276700
rect 302436 227050 302464 316006
rect 302424 227044 302476 227050
rect 302424 226986 302476 226992
rect 301504 18624 301556 18630
rect 301504 18566 301556 18572
rect 300860 11824 300912 11830
rect 300860 11766 300912 11772
rect 302896 6186 302924 336398
rect 302976 336320 303028 336326
rect 302976 336262 303028 336268
rect 302988 19990 303016 336262
rect 303080 333266 303108 336466
rect 303068 333260 303120 333266
rect 303068 333202 303120 333208
rect 303172 330546 303200 338014
rect 303160 330540 303212 330546
rect 303160 330482 303212 330488
rect 303724 267034 303752 338014
rect 303908 335354 303936 338014
rect 304276 336818 304304 338014
rect 304092 336790 304304 336818
rect 304092 336734 304120 336790
rect 304080 336728 304132 336734
rect 304644 336682 304672 338014
rect 304080 336670 304132 336676
rect 303816 335326 303936 335354
rect 304184 336654 304672 336682
rect 303816 319462 303844 335326
rect 303804 319456 303856 319462
rect 303804 319398 303856 319404
rect 304184 316034 304212 336654
rect 304264 335368 304316 335374
rect 304264 335310 304316 335316
rect 303908 316006 304212 316034
rect 303712 267028 303764 267034
rect 303712 266970 303764 266976
rect 303620 252068 303672 252074
rect 303620 252010 303672 252016
rect 302976 19984 303028 19990
rect 302976 19926 303028 19932
rect 303632 16574 303660 252010
rect 303908 251938 303936 316006
rect 303896 251932 303948 251938
rect 303896 251874 303948 251880
rect 303632 16546 303936 16574
rect 302884 6180 302936 6186
rect 302884 6122 302936 6128
rect 303160 5228 303212 5234
rect 303160 5170 303212 5176
rect 299664 5160 299716 5166
rect 299664 5102 299716 5108
rect 299480 2100 299532 2106
rect 299480 2042 299532 2048
rect 299676 480 299704 5102
rect 301964 4072 302016 4078
rect 301964 4014 302016 4020
rect 300768 2100 300820 2106
rect 300768 2042 300820 2048
rect 300780 480 300808 2042
rect 301976 480 302004 4014
rect 303172 480 303200 5170
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304276 7682 304304 335310
rect 305092 330540 305144 330546
rect 305092 330482 305144 330488
rect 305104 250578 305132 330482
rect 305196 318102 305224 338014
rect 305380 336530 305408 338014
rect 305368 336524 305420 336530
rect 305368 336466 305420 336472
rect 305644 335980 305696 335986
rect 305644 335922 305696 335928
rect 305276 326052 305328 326058
rect 305276 325994 305328 326000
rect 305184 318096 305236 318102
rect 305184 318038 305236 318044
rect 305092 250572 305144 250578
rect 305092 250514 305144 250520
rect 305288 240786 305316 325994
rect 305276 240780 305328 240786
rect 305276 240722 305328 240728
rect 304264 7676 304316 7682
rect 304264 7618 304316 7624
rect 305656 6254 305684 335922
rect 305748 330546 305776 338014
rect 305828 336388 305880 336394
rect 305828 336330 305880 336336
rect 305736 330540 305788 330546
rect 305736 330482 305788 330488
rect 305840 316034 305868 336330
rect 306116 326058 306144 338014
rect 306484 335354 306512 338014
rect 306852 335354 306880 338014
rect 307024 336252 307076 336258
rect 307024 336194 307076 336200
rect 306392 335326 306512 335354
rect 306668 335326 306880 335354
rect 306104 326052 306156 326058
rect 306104 325994 306156 326000
rect 306392 320890 306420 335326
rect 306668 330834 306696 335326
rect 306484 330806 306696 330834
rect 306380 320884 306432 320890
rect 306380 320826 306432 320832
rect 305748 316006 305868 316034
rect 305748 9110 305776 316006
rect 306484 247790 306512 330806
rect 306656 330540 306708 330546
rect 306656 330482 306708 330488
rect 306564 320884 306616 320890
rect 306564 320826 306616 320832
rect 306576 275398 306604 320826
rect 306564 275392 306616 275398
rect 306564 275334 306616 275340
rect 306472 247784 306524 247790
rect 306472 247726 306524 247732
rect 306668 17406 306696 330482
rect 307036 35222 307064 336194
rect 307220 335986 307248 338014
rect 307208 335980 307260 335986
rect 307208 335922 307260 335928
rect 307496 330546 307524 338014
rect 307864 335374 307892 338014
rect 307852 335368 307904 335374
rect 307852 335310 307904 335316
rect 307484 330540 307536 330546
rect 307484 330482 307536 330488
rect 308232 316034 308260 338014
rect 308600 335510 308628 338014
rect 309324 336728 309376 336734
rect 309324 336670 309376 336676
rect 308588 335504 308640 335510
rect 308588 335446 308640 335452
rect 309232 330540 309284 330546
rect 309232 330482 309284 330488
rect 307864 316006 308260 316034
rect 307864 44878 307892 316006
rect 307852 44872 307904 44878
rect 307852 44814 307904 44820
rect 307024 35216 307076 35222
rect 307024 35158 307076 35164
rect 309244 28286 309272 330482
rect 309336 46238 309364 336670
rect 309324 46232 309376 46238
rect 309324 46174 309376 46180
rect 309232 28280 309284 28286
rect 309232 28222 309284 28228
rect 309428 26926 309456 338150
rect 309520 338014 309580 338042
rect 309704 338014 309948 338042
rect 310072 338014 310316 338042
rect 309520 336734 309548 338014
rect 309508 336728 309560 336734
rect 309508 336670 309560 336676
rect 309704 336462 309732 338014
rect 309692 336456 309744 336462
rect 309692 336398 309744 336404
rect 310072 330546 310100 338014
rect 310670 337770 310698 338028
rect 310808 338014 311052 338042
rect 311176 338014 311420 338042
rect 311544 338014 311788 338042
rect 311912 338014 312156 338042
rect 312280 338014 312524 338042
rect 312648 338014 312892 338042
rect 313016 338014 313260 338042
rect 313384 338014 313628 338042
rect 313752 338014 313996 338042
rect 314120 338014 314364 338042
rect 310670 337742 310744 337770
rect 310060 330540 310112 330546
rect 310060 330482 310112 330488
rect 310612 330540 310664 330546
rect 310612 330482 310664 330488
rect 310624 29714 310652 330482
rect 310716 47598 310744 337742
rect 310808 336122 310836 338014
rect 310796 336116 310848 336122
rect 310796 336058 310848 336064
rect 311176 330546 311204 338014
rect 311164 330540 311216 330546
rect 311164 330482 311216 330488
rect 311544 316034 311572 338014
rect 311912 336190 311940 338014
rect 312280 336682 312308 338014
rect 312004 336654 312308 336682
rect 311900 336184 311952 336190
rect 311900 336126 311952 336132
rect 310808 316006 311572 316034
rect 310704 47592 310756 47598
rect 310704 47534 310756 47540
rect 310612 29708 310664 29714
rect 310612 29650 310664 29656
rect 310704 29640 310756 29646
rect 310704 29582 310756 29588
rect 309416 26920 309468 26926
rect 309416 26862 309468 26868
rect 307760 18624 307812 18630
rect 307760 18566 307812 18572
rect 306656 17400 306708 17406
rect 306656 17342 306708 17348
rect 306472 17264 306524 17270
rect 306472 17206 306524 17212
rect 305736 9104 305788 9110
rect 305736 9046 305788 9052
rect 305644 6248 305696 6254
rect 305644 6190 305696 6196
rect 305552 4140 305604 4146
rect 305552 4082 305604 4088
rect 305564 480 305592 4082
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306484 354 306512 17206
rect 307772 16574 307800 18566
rect 310716 16574 310744 29582
rect 310808 18698 310836 316006
rect 312004 31074 312032 336654
rect 312648 335354 312676 338014
rect 312096 335326 312676 335354
rect 312096 49026 312124 335326
rect 313016 316034 313044 338014
rect 313384 336394 313412 338014
rect 313372 336388 313424 336394
rect 313372 336330 313424 336336
rect 313372 330540 313424 330546
rect 313372 330482 313424 330488
rect 312188 316006 313044 316034
rect 312084 49020 312136 49026
rect 312084 48962 312136 48968
rect 311992 31068 312044 31074
rect 311992 31010 312044 31016
rect 312188 21418 312216 316006
rect 313384 22846 313412 330482
rect 313752 316034 313780 338014
rect 313924 335368 313976 335374
rect 313924 335310 313976 335316
rect 313476 316006 313780 316034
rect 313372 22840 313424 22846
rect 313372 22782 313424 22788
rect 312176 21412 312228 21418
rect 312176 21354 312228 21360
rect 310796 18692 310848 18698
rect 310796 18634 310848 18640
rect 313476 17338 313504 316006
rect 313464 17332 313516 17338
rect 313464 17274 313516 17280
rect 307772 16546 307984 16574
rect 310716 16546 311480 16574
rect 307956 480 307984 16546
rect 310244 7676 310296 7682
rect 310244 7618 310296 7624
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 7618
rect 311452 480 311480 16546
rect 313832 14544 313884 14550
rect 313832 14486 313884 14492
rect 312636 3324 312688 3330
rect 312636 3266 312688 3272
rect 312648 480 312676 3266
rect 313844 480 313872 14486
rect 313936 14482 313964 335310
rect 314120 330546 314148 338014
rect 314718 337770 314746 338028
rect 314856 338014 315100 338042
rect 315224 338014 315468 338042
rect 315592 338014 315836 338042
rect 316144 338014 316204 338042
rect 316328 338014 316572 338042
rect 316696 338014 316940 338042
rect 317064 338014 317308 338042
rect 317432 338014 317676 338042
rect 317800 338014 318044 338042
rect 318168 338014 318412 338042
rect 318536 338014 318780 338042
rect 318904 338014 319148 338042
rect 319272 338014 319424 338042
rect 319548 338014 319792 338042
rect 319916 338014 320160 338042
rect 320284 338014 320528 338042
rect 320652 338014 320896 338042
rect 321020 338014 321264 338042
rect 314718 337742 314792 337770
rect 314108 330540 314160 330546
rect 314108 330482 314160 330488
rect 314764 32434 314792 337742
rect 314856 336326 314884 338014
rect 314844 336320 314896 336326
rect 314844 336262 314896 336268
rect 315224 336054 315252 338014
rect 315304 336320 315356 336326
rect 315304 336262 315356 336268
rect 315212 336048 315264 336054
rect 315212 335990 315264 335996
rect 314844 330540 314896 330546
rect 314844 330482 314896 330488
rect 314752 32428 314804 32434
rect 314752 32370 314804 32376
rect 313924 14476 313976 14482
rect 313924 14418 313976 14424
rect 314856 10334 314884 330482
rect 314844 10328 314896 10334
rect 314844 10270 314896 10276
rect 315316 7614 315344 336262
rect 315592 330546 315620 338014
rect 315580 330540 315632 330546
rect 315580 330482 315632 330488
rect 316040 330472 316092 330478
rect 316040 330414 316092 330420
rect 315304 7608 315356 7614
rect 315304 7550 315356 7556
rect 316052 3466 316080 330414
rect 316144 25634 316172 338014
rect 316224 330540 316276 330546
rect 316224 330482 316276 330488
rect 316236 33794 316264 330482
rect 316328 180130 316356 338014
rect 316696 330546 316724 338014
rect 316684 330540 316736 330546
rect 316684 330482 316736 330488
rect 317064 330478 317092 338014
rect 317432 335374 317460 338014
rect 317420 335368 317472 335374
rect 317800 335354 317828 338014
rect 317420 335310 317472 335316
rect 317616 335326 317828 335354
rect 317052 330472 317104 330478
rect 317052 330414 317104 330420
rect 317512 330336 317564 330342
rect 317512 330278 317564 330284
rect 316316 180124 316368 180130
rect 316316 180066 316368 180072
rect 316224 33788 316276 33794
rect 316224 33730 316276 33736
rect 316132 25628 316184 25634
rect 316132 25570 316184 25576
rect 317524 13122 317552 330278
rect 317616 24206 317644 335326
rect 318168 316034 318196 338014
rect 318536 330342 318564 338014
rect 318800 330540 318852 330546
rect 318800 330482 318852 330488
rect 318524 330336 318576 330342
rect 318524 330278 318576 330284
rect 317708 316006 318196 316034
rect 317604 24200 317656 24206
rect 317604 24142 317656 24148
rect 317512 13116 317564 13122
rect 317512 13058 317564 13064
rect 317328 8968 317380 8974
rect 317328 8910 317380 8916
rect 316040 3460 316092 3466
rect 316040 3402 316092 3408
rect 315028 3256 315080 3262
rect 315028 3198 315080 3204
rect 315040 480 315068 3198
rect 316224 3188 316276 3194
rect 316224 3130 316276 3136
rect 316236 480 316264 3130
rect 317340 480 317368 8910
rect 317708 3534 317736 316006
rect 318812 3602 318840 330482
rect 318904 11762 318932 338014
rect 319272 330546 319300 338014
rect 319548 336682 319576 338014
rect 319364 336654 319576 336682
rect 319260 330540 319312 330546
rect 319260 330482 319312 330488
rect 318984 328228 319036 328234
rect 318984 328170 319036 328176
rect 318996 249218 319024 328170
rect 319364 316034 319392 336654
rect 319444 335844 319496 335850
rect 319444 335786 319496 335792
rect 319088 316006 319392 316034
rect 319088 274106 319116 316006
rect 319076 274100 319128 274106
rect 319076 274042 319128 274048
rect 318984 249212 319036 249218
rect 318984 249154 319036 249160
rect 319456 15910 319484 335786
rect 319916 328234 319944 338014
rect 320180 336048 320232 336054
rect 320180 335990 320232 335996
rect 319904 328228 319956 328234
rect 319904 328170 319956 328176
rect 319444 15904 319496 15910
rect 319444 15846 319496 15852
rect 318892 11756 318944 11762
rect 318892 11698 318944 11704
rect 318800 3596 318852 3602
rect 318800 3538 318852 3544
rect 317696 3528 317748 3534
rect 317696 3470 317748 3476
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 318524 3460 318576 3466
rect 318524 3402 318576 3408
rect 318536 480 318564 3402
rect 319732 480 319760 3470
rect 320192 490 320220 335990
rect 320284 3369 320312 338014
rect 320652 316034 320680 338014
rect 321020 335850 321048 338014
rect 321618 337770 321646 338028
rect 321756 338014 322000 338042
rect 322124 338014 322368 338042
rect 322492 338014 322736 338042
rect 321618 337742 321692 337770
rect 321008 335844 321060 335850
rect 321008 335786 321060 335792
rect 320824 335504 320876 335510
rect 320824 335446 320876 335452
rect 320376 316006 320680 316034
rect 320376 4894 320404 316006
rect 320836 253434 320864 335446
rect 321664 335238 321692 337742
rect 321652 335232 321704 335238
rect 321652 335174 321704 335180
rect 321652 326392 321704 326398
rect 321652 326334 321704 326340
rect 320824 253428 320876 253434
rect 320824 253370 320876 253376
rect 320364 4888 320416 4894
rect 320364 4830 320416 4836
rect 321664 3738 321692 326334
rect 321756 6322 321784 338014
rect 322124 336258 322152 338014
rect 322112 336252 322164 336258
rect 322112 336194 322164 336200
rect 322204 335708 322256 335714
rect 322204 335650 322256 335656
rect 321836 335232 321888 335238
rect 321836 335174 321888 335180
rect 321744 6316 321796 6322
rect 321744 6258 321796 6264
rect 321652 3732 321704 3738
rect 321652 3674 321704 3680
rect 321848 3670 321876 335174
rect 322216 279682 322244 335650
rect 322492 326398 322520 338014
rect 323090 337770 323118 338028
rect 323228 338014 323472 338042
rect 323596 338014 323840 338042
rect 323964 338014 324208 338042
rect 324332 338014 324576 338042
rect 324700 338014 324944 338042
rect 325068 338014 325312 338042
rect 325436 338014 325680 338042
rect 325896 338014 326048 338042
rect 326172 338014 326416 338042
rect 326540 338014 326784 338042
rect 323090 337742 323164 337770
rect 323032 326460 323084 326466
rect 323032 326402 323084 326408
rect 322480 326392 322532 326398
rect 322480 326334 322532 326340
rect 322940 326392 322992 326398
rect 322940 326334 322992 326340
rect 322204 279676 322256 279682
rect 322204 279618 322256 279624
rect 322952 3806 322980 326334
rect 323044 5030 323072 326402
rect 323032 5024 323084 5030
rect 323032 4966 323084 4972
rect 323136 4962 323164 337742
rect 323228 284986 323256 338014
rect 323596 326398 323624 338014
rect 323964 326466 323992 338014
rect 324332 336326 324360 338014
rect 324700 336682 324728 338014
rect 324424 336654 324728 336682
rect 324320 336320 324372 336326
rect 324320 336262 324372 336268
rect 324320 336184 324372 336190
rect 324320 336126 324372 336132
rect 323952 326460 324004 326466
rect 323952 326402 324004 326408
rect 323584 326392 323636 326398
rect 323584 326334 323636 326340
rect 323216 284980 323268 284986
rect 323216 284922 323268 284928
rect 323124 4956 323176 4962
rect 323124 4898 323176 4904
rect 322940 3800 322992 3806
rect 322940 3742 322992 3748
rect 323308 3732 323360 3738
rect 323308 3674 323360 3680
rect 321836 3664 321888 3670
rect 321836 3606 321888 3612
rect 322112 3596 322164 3602
rect 322112 3538 322164 3544
rect 320270 3360 320326 3369
rect 320270 3295 320326 3304
rect 306718 354 306830 480
rect 306484 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320192 462 320496 490
rect 322124 480 322152 3538
rect 323320 480 323348 3674
rect 324332 3482 324360 336126
rect 324424 3874 324452 336654
rect 325068 335354 325096 338014
rect 324516 335326 325096 335354
rect 324516 4826 324544 335326
rect 325436 316034 325464 338014
rect 325896 328454 325924 338014
rect 326172 335354 326200 338014
rect 326540 335714 326568 338014
rect 327138 337770 327166 338028
rect 327368 338014 327520 338042
rect 327644 338014 327888 338042
rect 328012 338014 328256 338042
rect 328564 338014 328624 338042
rect 328748 338014 328992 338042
rect 329116 338014 329360 338042
rect 329484 338014 329728 338042
rect 330036 338014 330096 338042
rect 330220 338014 330464 338042
rect 330588 338014 330832 338042
rect 330956 338014 331108 338042
rect 331416 338014 331476 338042
rect 331600 338014 331844 338042
rect 331968 338014 332212 338042
rect 332336 338014 332580 338042
rect 332796 338014 332948 338042
rect 333072 338014 333316 338042
rect 333440 338014 333684 338042
rect 333992 338014 334052 338042
rect 334176 338014 334420 338042
rect 334544 338014 334788 338042
rect 334912 338014 335156 338042
rect 327138 337742 327212 337770
rect 327080 336116 327132 336122
rect 327080 336058 327132 336064
rect 326528 335708 326580 335714
rect 326528 335650 326580 335656
rect 325804 328426 325924 328454
rect 325988 335326 326200 335354
rect 325804 323762 325832 328426
rect 325804 323734 325924 323762
rect 325792 323604 325844 323610
rect 325792 323546 325844 323552
rect 324608 316006 325464 316034
rect 324608 261594 324636 316006
rect 324596 261588 324648 261594
rect 324596 261530 324648 261536
rect 325804 5098 325832 323546
rect 325792 5092 325844 5098
rect 325792 5034 325844 5040
rect 324504 4820 324556 4826
rect 324504 4762 324556 4768
rect 325896 3942 325924 323734
rect 325988 323610 326016 335326
rect 325976 323604 326028 323610
rect 325976 323546 326028 323552
rect 325884 3936 325936 3942
rect 325884 3878 325936 3884
rect 324412 3868 324464 3874
rect 324412 3810 324464 3816
rect 326804 3800 326856 3806
rect 326804 3742 326856 3748
rect 325608 3664 325660 3670
rect 325608 3606 325660 3612
rect 324332 3454 324452 3482
rect 324424 480 324452 3454
rect 325620 480 325648 3606
rect 326816 480 326844 3742
rect 327092 3482 327120 336058
rect 327184 4010 327212 337742
rect 327264 326392 327316 326398
rect 327264 326334 327316 326340
rect 327276 4078 327304 326334
rect 327368 5166 327396 338014
rect 327644 335510 327672 338014
rect 327632 335504 327684 335510
rect 327632 335446 327684 335452
rect 328012 326398 328040 338014
rect 328460 326460 328512 326466
rect 328460 326402 328512 326408
rect 328000 326392 328052 326398
rect 328000 326334 328052 326340
rect 327356 5160 327408 5166
rect 327356 5102 327408 5108
rect 328472 4146 328500 326402
rect 328564 5234 328592 338014
rect 328644 326392 328696 326398
rect 328644 326334 328696 326340
rect 328656 17270 328684 326334
rect 328748 252074 328776 338014
rect 329116 326466 329144 338014
rect 329104 326460 329156 326466
rect 329104 326402 329156 326408
rect 329484 326398 329512 338014
rect 329472 326392 329524 326398
rect 329472 326334 329524 326340
rect 329932 326392 329984 326398
rect 329932 326334 329984 326340
rect 329840 321632 329892 321638
rect 329840 321574 329892 321580
rect 328736 252068 328788 252074
rect 328736 252010 328788 252016
rect 328644 17264 328696 17270
rect 328644 17206 328696 17212
rect 328552 5228 328604 5234
rect 328552 5170 328604 5176
rect 328460 4140 328512 4146
rect 328460 4082 328512 4088
rect 327264 4072 327316 4078
rect 327264 4014 327316 4020
rect 327172 4004 327224 4010
rect 327172 3946 327224 3952
rect 329012 3868 329064 3874
rect 329012 3810 329064 3816
rect 329024 3602 329052 3810
rect 329012 3596 329064 3602
rect 329012 3538 329064 3544
rect 327092 3454 328040 3482
rect 328012 480 328040 3454
rect 329852 3398 329880 321574
rect 329944 7682 329972 326334
rect 330036 18630 330064 338014
rect 330220 321638 330248 338014
rect 330588 326398 330616 338014
rect 330576 326392 330628 326398
rect 330576 326334 330628 326340
rect 330208 321632 330260 321638
rect 330208 321574 330260 321580
rect 330956 316034 330984 338014
rect 331220 330540 331272 330546
rect 331220 330482 331272 330488
rect 330128 316006 330984 316034
rect 330128 29646 330156 316006
rect 330116 29640 330168 29646
rect 330116 29582 330168 29588
rect 330024 18624 330076 18630
rect 330024 18566 330076 18572
rect 329932 7676 329984 7682
rect 329932 7618 329984 7624
rect 330392 4004 330444 4010
rect 330392 3946 330444 3952
rect 329840 3392 329892 3398
rect 329840 3334 329892 3340
rect 329196 3052 329248 3058
rect 329196 2994 329248 3000
rect 329208 480 329236 2994
rect 330404 480 330432 3946
rect 331232 3262 331260 330482
rect 331312 330472 331364 330478
rect 331312 330414 331364 330420
rect 331220 3256 331272 3262
rect 331220 3198 331272 3204
rect 331324 3194 331352 330414
rect 331416 3330 331444 338014
rect 331600 316034 331628 338014
rect 331968 330546 331996 338014
rect 331956 330540 332008 330546
rect 331956 330482 332008 330488
rect 332336 330478 332364 338014
rect 332600 330540 332652 330546
rect 332600 330482 332652 330488
rect 332324 330472 332376 330478
rect 332324 330414 332376 330420
rect 331508 316006 331628 316034
rect 331508 14550 331536 316006
rect 331496 14544 331548 14550
rect 331496 14486 331548 14492
rect 332612 3602 332640 330482
rect 332692 327548 332744 327554
rect 332692 327490 332744 327496
rect 332704 6914 332732 327490
rect 332796 8974 332824 338014
rect 333072 327554 333100 338014
rect 333244 335368 333296 335374
rect 333244 335310 333296 335316
rect 333060 327548 333112 327554
rect 333060 327490 333112 327496
rect 332784 8968 332836 8974
rect 332784 8910 332836 8916
rect 332704 6886 332824 6914
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 332600 3596 332652 3602
rect 332600 3538 332652 3544
rect 331588 3528 331640 3534
rect 331588 3470 331640 3476
rect 331404 3324 331456 3330
rect 331404 3266 331456 3272
rect 331312 3188 331364 3194
rect 331312 3130 331364 3136
rect 331600 480 331628 3470
rect 332704 480 332732 4014
rect 332796 3466 332824 6886
rect 333256 3534 333284 335310
rect 333440 330546 333468 338014
rect 333992 336054 334020 338014
rect 333980 336048 334032 336054
rect 333980 335990 334032 335996
rect 333428 330540 333480 330546
rect 333428 330482 333480 330488
rect 334072 330540 334124 330546
rect 334072 330482 334124 330488
rect 333888 4140 333940 4146
rect 333888 4082 333940 4088
rect 333244 3528 333296 3534
rect 333244 3470 333296 3476
rect 332784 3460 332836 3466
rect 332784 3402 332836 3408
rect 333900 480 333928 4082
rect 334084 3738 334112 330482
rect 334176 3874 334204 338014
rect 334348 336320 334400 336326
rect 334348 336262 334400 336268
rect 334360 16574 334388 336262
rect 334544 330546 334572 338014
rect 334912 336190 334940 338014
rect 335510 337770 335538 338028
rect 335648 338014 335892 338042
rect 336016 338014 336260 338042
rect 336384 338014 336628 338042
rect 336936 338014 336996 338042
rect 337120 338014 337364 338042
rect 337488 338014 337732 338042
rect 337856 338014 338100 338042
rect 338224 338014 338468 338042
rect 338592 338014 338836 338042
rect 338960 338014 339204 338042
rect 335510 337742 335584 337770
rect 335452 336728 335504 336734
rect 335452 336670 335504 336676
rect 334900 336184 334952 336190
rect 334900 336126 334952 336132
rect 334532 330540 334584 330546
rect 334532 330482 334584 330488
rect 334360 16546 334664 16574
rect 334164 3868 334216 3874
rect 334164 3810 334216 3816
rect 334072 3732 334124 3738
rect 334072 3674 334124 3680
rect 320468 354 320496 462
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335464 3806 335492 336670
rect 335452 3800 335504 3806
rect 335452 3742 335504 3748
rect 335556 3670 335584 337742
rect 335648 336734 335676 338014
rect 335636 336728 335688 336734
rect 335636 336670 335688 336676
rect 336016 336122 336044 338014
rect 336004 336116 336056 336122
rect 336004 336058 336056 336064
rect 336384 316034 336412 338014
rect 336832 330540 336884 330546
rect 336832 330482 336884 330488
rect 335648 316006 336412 316034
rect 335544 3664 335596 3670
rect 335544 3606 335596 3612
rect 335648 3058 335676 316006
rect 336844 4146 336872 330482
rect 336832 4140 336884 4146
rect 336832 4082 336884 4088
rect 336936 4010 336964 338014
rect 337120 335374 337148 338014
rect 337108 335368 337160 335374
rect 337108 335310 337160 335316
rect 337488 316034 337516 338014
rect 337856 330546 337884 338014
rect 338224 336326 338252 338014
rect 338212 336320 338264 336326
rect 338212 336262 338264 336268
rect 338592 335354 338620 338014
rect 338316 335326 338620 335354
rect 337844 330540 337896 330546
rect 337844 330482 337896 330488
rect 338316 316034 338344 335326
rect 338960 316034 338988 338014
rect 339558 337770 339586 338028
rect 339696 338014 339940 338042
rect 340064 338014 340308 338042
rect 340676 338014 340828 338042
rect 339558 337742 339632 337770
rect 339500 336252 339552 336258
rect 339500 336194 339552 336200
rect 337120 316006 337516 316034
rect 338224 316006 338344 316034
rect 338408 316006 338988 316034
rect 337120 4078 337148 316006
rect 337108 4072 337160 4078
rect 337108 4014 337160 4020
rect 336924 4004 336976 4010
rect 336924 3946 336976 3952
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 336280 3188 336332 3194
rect 336280 3130 336332 3136
rect 335636 3052 335688 3058
rect 335636 2994 335688 3000
rect 336292 480 336320 3130
rect 337488 480 337516 3470
rect 338224 3194 338252 316006
rect 338408 3534 338436 316006
rect 338396 3528 338448 3534
rect 338396 3470 338448 3476
rect 338672 3528 338724 3534
rect 338672 3470 338724 3476
rect 338212 3188 338264 3194
rect 338212 3130 338264 3136
rect 338684 480 338712 3470
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 336194
rect 339604 3534 339632 337742
rect 339696 336258 339724 338014
rect 339684 336252 339736 336258
rect 339684 336194 339736 336200
rect 340064 316034 340092 338014
rect 340800 336598 340828 338014
rect 340984 338014 341044 338042
rect 341168 338014 341412 338042
rect 341536 338014 341780 338042
rect 341904 338014 342148 338042
rect 342364 338014 342516 338042
rect 342640 338014 342884 338042
rect 343008 338014 343160 338042
rect 343284 338014 343528 338042
rect 343836 338014 343896 338042
rect 344020 338014 344264 338042
rect 344388 338014 344632 338042
rect 344940 338014 345000 338042
rect 345124 338014 345368 338042
rect 340788 336592 340840 336598
rect 340788 336534 340840 336540
rect 340984 335714 341012 338014
rect 340972 335708 341024 335714
rect 340972 335650 341024 335656
rect 341168 330528 341196 338014
rect 341536 336682 341564 338014
rect 341076 330500 341196 330528
rect 341260 336654 341564 336682
rect 340972 329860 341024 329866
rect 340972 329802 341024 329808
rect 339696 316006 340092 316034
rect 339696 3534 339724 316006
rect 340984 6914 341012 329802
rect 340892 6886 341012 6914
rect 340892 4078 340920 6886
rect 340880 4072 340932 4078
rect 340880 4014 340932 4020
rect 339592 3528 339644 3534
rect 339592 3470 339644 3476
rect 339684 3528 339736 3534
rect 339684 3470 339736 3476
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 340984 480 341012 3470
rect 341076 3398 341104 330500
rect 341260 316034 341288 336654
rect 341340 336592 341392 336598
rect 341340 336534 341392 336540
rect 341168 316006 341288 316034
rect 341064 3392 341116 3398
rect 341064 3334 341116 3340
rect 341168 2922 341196 316006
rect 341352 16574 341380 336534
rect 341904 329866 341932 338014
rect 342260 335708 342312 335714
rect 342260 335650 342312 335656
rect 341892 329860 341944 329866
rect 341892 329802 341944 329808
rect 341352 16546 342208 16574
rect 341156 2916 341208 2922
rect 341156 2858 341208 2864
rect 342180 480 342208 16546
rect 342272 762 342300 335650
rect 342364 3806 342392 338014
rect 342536 330540 342588 330546
rect 342536 330482 342588 330488
rect 342444 330472 342496 330478
rect 342444 330414 342496 330420
rect 342352 3800 342404 3806
rect 342352 3742 342404 3748
rect 342456 3602 342484 330414
rect 342548 3738 342576 330482
rect 342640 3874 342668 338014
rect 343008 330546 343036 338014
rect 342996 330540 343048 330546
rect 342996 330482 343048 330488
rect 343284 330478 343312 338014
rect 343836 336326 343864 338014
rect 343824 336320 343876 336326
rect 343824 336262 343876 336268
rect 344020 335354 344048 338014
rect 343652 335326 344048 335354
rect 343272 330472 343324 330478
rect 343272 330414 343324 330420
rect 342628 3868 342680 3874
rect 342628 3810 342680 3816
rect 342536 3732 342588 3738
rect 342536 3674 342588 3680
rect 342444 3596 342496 3602
rect 342444 3538 342496 3544
rect 343652 3534 343680 335326
rect 344388 316034 344416 338014
rect 344940 336054 344968 338014
rect 344928 336048 344980 336054
rect 344928 335990 344980 335996
rect 345020 330540 345072 330546
rect 345020 330482 345072 330488
rect 343744 316006 344416 316034
rect 343640 3528 343692 3534
rect 343640 3470 343692 3476
rect 343744 3466 343772 316006
rect 345032 6254 345060 330482
rect 345124 10402 345152 338014
rect 345722 337770 345750 338028
rect 345860 338014 346104 338042
rect 346472 338014 346624 338042
rect 345722 337742 345796 337770
rect 345768 336326 345796 337742
rect 345664 336320 345716 336326
rect 345664 336262 345716 336268
rect 345756 336320 345808 336326
rect 345756 336262 345808 336268
rect 345112 10396 345164 10402
rect 345112 10338 345164 10344
rect 345020 6248 345072 6254
rect 345020 6190 345072 6196
rect 345676 4214 345704 336262
rect 345860 330546 345888 338014
rect 346400 336728 346452 336734
rect 346400 336670 346452 336676
rect 345848 330540 345900 330546
rect 345848 330482 345900 330488
rect 345664 4208 345716 4214
rect 345664 4150 345716 4156
rect 346412 3670 346440 336670
rect 346492 327820 346544 327826
rect 346492 327762 346544 327768
rect 346504 6186 346532 327762
rect 346596 17270 346624 338014
rect 346688 338014 346840 338042
rect 347208 338014 347360 338042
rect 346688 336734 346716 338014
rect 346676 336728 346728 336734
rect 346676 336670 346728 336676
rect 347332 336258 347360 338014
rect 347424 338014 347576 338042
rect 347320 336252 347372 336258
rect 347320 336194 347372 336200
rect 347424 327826 347452 338014
rect 347930 337770 347958 338028
rect 348068 338014 348312 338042
rect 348620 338014 348680 338042
rect 348804 338014 349048 338042
rect 349172 338014 349416 338042
rect 349540 338014 349784 338042
rect 350092 338014 350152 338042
rect 350276 338014 350520 338042
rect 350828 338014 350888 338042
rect 351012 338014 351256 338042
rect 351380 338014 351624 338042
rect 351932 338014 351992 338042
rect 352116 338014 352360 338042
rect 352484 338014 352728 338042
rect 352852 338014 353096 338042
rect 353312 338014 353464 338042
rect 353772 338014 353832 338042
rect 353956 338014 354200 338042
rect 354324 338014 354568 338042
rect 347930 337742 348004 337770
rect 347976 330818 348004 337742
rect 347964 330812 348016 330818
rect 347964 330754 348016 330760
rect 348068 330698 348096 338014
rect 348620 336190 348648 338014
rect 348608 336184 348660 336190
rect 348608 336126 348660 336132
rect 347792 330670 348096 330698
rect 347412 327820 347464 327826
rect 347412 327762 347464 327768
rect 346584 17264 346636 17270
rect 346584 17206 346636 17212
rect 347792 7682 347820 330670
rect 347964 330608 348016 330614
rect 347964 330550 348016 330556
rect 347872 330540 347924 330546
rect 347872 330482 347924 330488
rect 347884 18630 347912 330482
rect 347976 51746 348004 330550
rect 348804 330546 348832 338014
rect 348792 330540 348844 330546
rect 348792 330482 348844 330488
rect 347964 51740 348016 51746
rect 347964 51682 348016 51688
rect 347872 18624 347924 18630
rect 347872 18566 347924 18572
rect 349172 9042 349200 338014
rect 349540 335354 349568 338014
rect 350092 336530 350120 338014
rect 350080 336524 350132 336530
rect 350080 336466 350132 336472
rect 349264 335326 349568 335354
rect 349264 10334 349292 335326
rect 350276 316034 350304 338014
rect 350828 336122 350856 338014
rect 350816 336116 350868 336122
rect 350816 336058 350868 336064
rect 350540 326392 350592 326398
rect 350540 326334 350592 326340
rect 349356 316006 350304 316034
rect 349356 11830 349384 316006
rect 350552 13122 350580 326334
rect 351012 316034 351040 338014
rect 351184 336048 351236 336054
rect 351184 335990 351236 335996
rect 350644 316006 351040 316034
rect 350644 26926 350672 316006
rect 350632 26920 350684 26926
rect 350632 26862 350684 26868
rect 350540 13116 350592 13122
rect 350540 13058 350592 13064
rect 349344 11824 349396 11830
rect 349344 11766 349396 11772
rect 349252 10328 349304 10334
rect 349252 10270 349304 10276
rect 349160 9036 349212 9042
rect 349160 8978 349212 8984
rect 347780 7676 347832 7682
rect 347780 7618 347832 7624
rect 346492 6180 346544 6186
rect 346492 6122 346544 6128
rect 351196 4894 351224 335990
rect 351380 326398 351408 338014
rect 351932 336054 351960 338014
rect 351920 336048 351972 336054
rect 351920 335990 351972 335996
rect 352116 335866 352144 338014
rect 351932 335838 352144 335866
rect 351368 326392 351420 326398
rect 351368 326334 351420 326340
rect 351932 7614 351960 335838
rect 352484 335354 352512 338014
rect 352024 335326 352512 335354
rect 352024 14482 352052 335326
rect 352852 316034 352880 338014
rect 352116 316006 352880 316034
rect 352116 21418 352144 316006
rect 352104 21412 352156 21418
rect 352104 21354 352156 21360
rect 352012 14476 352064 14482
rect 352012 14418 352064 14424
rect 353312 8974 353340 338014
rect 353772 336462 353800 338014
rect 353760 336456 353812 336462
rect 353760 336398 353812 336404
rect 353956 335354 353984 338014
rect 353404 335326 353984 335354
rect 353404 47598 353432 335326
rect 354324 316034 354352 338014
rect 354922 337770 354950 338028
rect 355060 338014 355212 338042
rect 355336 338014 355580 338042
rect 355704 338014 355948 338042
rect 356256 338014 356316 338042
rect 356440 338014 356684 338042
rect 356808 338014 357052 338042
rect 357176 338014 357420 338042
rect 357544 338014 357788 338042
rect 354922 337742 354996 337770
rect 354968 326534 354996 337742
rect 354956 326528 355008 326534
rect 354956 326470 355008 326476
rect 354680 326460 354732 326466
rect 354680 326402 354732 326408
rect 353496 316006 354352 316034
rect 353496 246362 353524 316006
rect 353484 246356 353536 246362
rect 353484 246298 353536 246304
rect 353392 47592 353444 47598
rect 353392 47534 353444 47540
rect 353300 8968 353352 8974
rect 353300 8910 353352 8916
rect 351920 7608 351972 7614
rect 351920 7550 351972 7556
rect 351184 4888 351236 4894
rect 351184 4830 351236 4836
rect 354692 4826 354720 326402
rect 354772 326392 354824 326398
rect 354772 326334 354824 326340
rect 354784 29646 354812 326334
rect 355060 323626 355088 338014
rect 355140 326528 355192 326534
rect 355140 326470 355192 326476
rect 354876 323598 355088 323626
rect 354876 261526 354904 323598
rect 355152 318794 355180 326470
rect 355336 326398 355364 338014
rect 355704 326466 355732 338014
rect 356256 326466 356284 338014
rect 356440 335354 356468 338014
rect 356348 335326 356468 335354
rect 355692 326460 355744 326466
rect 355692 326402 355744 326408
rect 356244 326460 356296 326466
rect 356244 326402 356296 326408
rect 355324 326392 355376 326398
rect 355324 326334 355376 326340
rect 356060 326392 356112 326398
rect 356060 326334 356112 326340
rect 354968 318766 355180 318794
rect 354968 286414 354996 318766
rect 354956 286408 355008 286414
rect 354956 286350 355008 286356
rect 354864 261520 354916 261526
rect 354864 261462 354916 261468
rect 354772 29640 354824 29646
rect 354772 29582 354824 29588
rect 356072 22778 356100 326334
rect 356348 323626 356376 335326
rect 356428 326460 356480 326466
rect 356428 326402 356480 326408
rect 356164 323598 356376 323626
rect 356164 28422 356192 323598
rect 356440 318794 356468 326402
rect 356256 318766 356468 318794
rect 356256 260166 356284 318766
rect 356808 316034 356836 338014
rect 357176 326398 357204 338014
rect 357440 336320 357492 336326
rect 357440 336262 357492 336268
rect 357164 326392 357216 326398
rect 357164 326334 357216 326340
rect 356348 316006 356836 316034
rect 356348 285054 356376 316006
rect 356336 285048 356388 285054
rect 356336 284990 356388 284996
rect 356244 260160 356296 260166
rect 356244 260102 356296 260108
rect 356152 28416 356204 28422
rect 356152 28358 356204 28364
rect 356060 22772 356112 22778
rect 356060 22714 356112 22720
rect 356336 4888 356388 4894
rect 356336 4830 356388 4836
rect 354680 4820 354732 4826
rect 354680 4762 354732 4768
rect 352840 4208 352892 4214
rect 352840 4150 352892 4156
rect 346952 4072 347004 4078
rect 346952 4014 347004 4020
rect 346400 3664 346452 3670
rect 346400 3606 346452 3612
rect 343732 3460 343784 3466
rect 343732 3402 343784 3408
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 342272 734 342944 762
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 734
rect 344572 480 344600 3334
rect 345756 2916 345808 2922
rect 345756 2858 345808 2864
rect 345768 480 345796 2858
rect 346964 480 346992 4014
rect 349252 3868 349304 3874
rect 349252 3810 349304 3816
rect 348056 3800 348108 3806
rect 348056 3742 348108 3748
rect 348068 480 348096 3742
rect 349264 480 349292 3810
rect 350448 3732 350500 3738
rect 350448 3674 350500 3680
rect 350460 480 350488 3674
rect 351644 3596 351696 3602
rect 351644 3538 351696 3544
rect 351656 480 351684 3538
rect 352852 480 352880 4150
rect 354036 3528 354088 3534
rect 354036 3470 354088 3476
rect 354048 480 354076 3470
rect 355232 3460 355284 3466
rect 355232 3402 355284 3408
rect 355244 480 355272 3402
rect 356348 480 356376 4830
rect 357452 3534 357480 336262
rect 357544 32434 357572 338014
rect 358142 337770 358170 338028
rect 358280 338014 358524 338042
rect 358892 338014 359044 338042
rect 358142 337742 358216 337770
rect 358084 336524 358136 336530
rect 358084 336466 358136 336472
rect 357624 322652 357676 322658
rect 357624 322594 357676 322600
rect 357636 256018 357664 322594
rect 357624 256012 357676 256018
rect 357624 255954 357676 255960
rect 357532 32428 357584 32434
rect 357532 32370 357584 32376
rect 358096 25566 358124 336466
rect 358188 336394 358216 337742
rect 358176 336388 358228 336394
rect 358176 336330 358228 336336
rect 358280 322658 358308 338014
rect 359016 331214 359044 338014
rect 358924 331186 359044 331214
rect 359108 338014 359260 338042
rect 359384 338014 359628 338042
rect 359752 338014 359996 338042
rect 360304 338014 360364 338042
rect 360488 338014 360732 338042
rect 360856 338014 361100 338042
rect 361224 338014 361468 338042
rect 361776 338014 361836 338042
rect 361960 338014 362204 338042
rect 362572 338014 362816 338042
rect 358924 323626 358952 331186
rect 358924 323598 359044 323626
rect 358912 323264 358964 323270
rect 358912 323206 358964 323212
rect 358268 322652 358320 322658
rect 358268 322594 358320 322600
rect 358820 322584 358872 322590
rect 358820 322526 358872 322532
rect 358084 25560 358136 25566
rect 358084 25502 358136 25508
rect 358832 15910 358860 322526
rect 358924 31074 358952 323206
rect 359016 254590 359044 323598
rect 359108 322590 359136 338014
rect 359096 322584 359148 322590
rect 359096 322526 359148 322532
rect 359384 316034 359412 338014
rect 359464 336184 359516 336190
rect 359464 336126 359516 336132
rect 359476 335986 359504 336126
rect 359464 335980 359516 335986
rect 359464 335922 359516 335928
rect 359752 323270 359780 338014
rect 360200 330540 360252 330546
rect 360200 330482 360252 330488
rect 359740 323264 359792 323270
rect 359740 323206 359792 323212
rect 359108 316006 359412 316034
rect 359108 272542 359136 316006
rect 359096 272536 359148 272542
rect 359096 272478 359148 272484
rect 359004 254584 359056 254590
rect 359004 254526 359056 254532
rect 358912 31068 358964 31074
rect 358912 31010 358964 31016
rect 358820 15904 358872 15910
rect 358820 15846 358872 15852
rect 357532 10396 357584 10402
rect 357532 10338 357584 10344
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 357544 480 357572 10338
rect 359924 6248 359976 6254
rect 359924 6190 359976 6196
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 358740 480 358768 3470
rect 359936 480 359964 6190
rect 360212 3602 360240 330482
rect 360304 17406 360332 338014
rect 360488 335354 360516 338014
rect 360396 335326 360516 335354
rect 360396 24138 360424 335326
rect 360856 330546 360884 338014
rect 360844 330540 360896 330546
rect 360844 330482 360896 330488
rect 361224 316034 361252 338014
rect 361776 335510 361804 338014
rect 361764 335504 361816 335510
rect 361764 335446 361816 335452
rect 361960 316034 361988 338014
rect 362788 336326 362816 338014
rect 362880 338014 362940 338042
rect 363064 338014 363308 338042
rect 363432 338014 363676 338042
rect 363800 338014 364044 338042
rect 364352 338014 364412 338042
rect 364628 338014 364780 338042
rect 364904 338014 365148 338042
rect 365272 338014 365516 338042
rect 362880 336530 362908 338014
rect 362868 336524 362920 336530
rect 362868 336466 362920 336472
rect 362776 336320 362828 336326
rect 362776 336262 362828 336268
rect 362960 336252 363012 336258
rect 362960 336194 363012 336200
rect 360488 316006 361252 316034
rect 361592 316006 361988 316034
rect 360488 283694 360516 316006
rect 360476 283688 360528 283694
rect 360476 283630 360528 283636
rect 360384 24132 360436 24138
rect 360384 24074 360436 24080
rect 360292 17400 360344 17406
rect 360292 17342 360344 17348
rect 360292 17264 360344 17270
rect 360292 17206 360344 17212
rect 360304 16574 360332 17206
rect 360304 16546 361160 16574
rect 360200 3596 360252 3602
rect 360200 3538 360252 3544
rect 361132 480 361160 16546
rect 361592 3466 361620 316006
rect 362972 6914 363000 336194
rect 363064 13190 363092 338014
rect 363432 335354 363460 338014
rect 363156 335326 363460 335354
rect 363156 282266 363184 335326
rect 363800 324970 363828 338014
rect 363788 324964 363840 324970
rect 363788 324906 363840 324912
rect 363144 282260 363196 282266
rect 363144 282202 363196 282208
rect 363052 13184 363104 13190
rect 363052 13126 363104 13132
rect 362972 6886 363552 6914
rect 362316 3664 362368 3670
rect 362316 3606 362368 3612
rect 361580 3460 361632 3466
rect 361580 3402 361632 3408
rect 362328 480 362356 3606
rect 363524 480 363552 6886
rect 364352 3262 364380 338014
rect 364432 330540 364484 330546
rect 364432 330482 364484 330488
rect 364444 3330 364472 330482
rect 364628 326398 364656 338014
rect 364616 326392 364668 326398
rect 364616 326334 364668 326340
rect 364904 321026 364932 338014
rect 364984 335504 365036 335510
rect 364984 335446 365036 335452
rect 364892 321020 364944 321026
rect 364892 320962 364944 320968
rect 364996 250510 365024 335446
rect 365272 330546 365300 338014
rect 365870 337770 365898 338028
rect 366238 337770 366266 338028
rect 366376 338014 366620 338042
rect 366744 338014 366988 338042
rect 367264 338014 367416 338042
rect 365870 337742 365944 337770
rect 366238 337742 366312 337770
rect 365260 330540 365312 330546
rect 365260 330482 365312 330488
rect 365812 329588 365864 329594
rect 365812 329530 365864 329536
rect 365720 327684 365772 327690
rect 365720 327626 365772 327632
rect 364984 250504 365036 250510
rect 364984 250446 365036 250452
rect 364616 6180 364668 6186
rect 364616 6122 364668 6128
rect 364432 3324 364484 3330
rect 364432 3266 364484 3272
rect 364340 3256 364392 3262
rect 364340 3198 364392 3204
rect 364628 480 364656 6122
rect 365732 3398 365760 327626
rect 365824 280906 365852 329530
rect 365916 298790 365944 337742
rect 366180 335980 366232 335986
rect 366180 335922 366232 335928
rect 366192 325694 366220 335922
rect 366284 330614 366312 337742
rect 366272 330608 366324 330614
rect 366272 330550 366324 330556
rect 366376 327690 366404 338014
rect 366744 329594 366772 338014
rect 367100 336728 367152 336734
rect 367100 336670 367152 336676
rect 366732 329588 366784 329594
rect 366732 329530 366784 329536
rect 366364 327684 366416 327690
rect 366364 327626 366416 327632
rect 366192 325666 366404 325694
rect 365904 298784 365956 298790
rect 365904 298726 365956 298732
rect 365812 280900 365864 280906
rect 365812 280842 365864 280848
rect 365812 51740 365864 51746
rect 365812 51682 365864 51688
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 51682
rect 366376 5574 366404 325666
rect 367008 7676 367060 7682
rect 367008 7618 367060 7624
rect 366364 5568 366416 5574
rect 366364 5510 366416 5516
rect 367020 480 367048 7618
rect 367112 4146 367140 336670
rect 367192 336660 367244 336666
rect 367192 336602 367244 336608
rect 367204 6526 367232 336602
rect 367284 330540 367336 330546
rect 367284 330482 367336 330488
rect 367296 258738 367324 330482
rect 367388 319530 367416 338014
rect 367480 338014 367632 338042
rect 367756 338014 368000 338042
rect 368124 338014 368368 338042
rect 368492 338014 368736 338042
rect 368860 338014 369104 338042
rect 369228 338014 369472 338042
rect 369596 338014 369840 338042
rect 369964 338014 370208 338042
rect 370332 338014 370576 338042
rect 370700 338014 370944 338042
rect 367480 336734 367508 338014
rect 367468 336728 367520 336734
rect 367468 336670 367520 336676
rect 367756 336666 367784 338014
rect 367744 336660 367796 336666
rect 367744 336602 367796 336608
rect 368124 330546 368152 338014
rect 368112 330540 368164 330546
rect 368112 330482 368164 330488
rect 367376 319524 367428 319530
rect 367376 319466 367428 319472
rect 367284 258732 367336 258738
rect 367284 258674 367336 258680
rect 367192 6520 367244 6526
rect 367192 6462 367244 6468
rect 368204 5568 368256 5574
rect 368204 5510 368256 5516
rect 367100 4140 367152 4146
rect 367100 4082 367152 4088
rect 368216 480 368244 5510
rect 368492 4078 368520 338014
rect 368860 335354 368888 338014
rect 368676 335326 368888 335354
rect 368572 330540 368624 330546
rect 368572 330482 368624 330488
rect 368480 4072 368532 4078
rect 368480 4014 368532 4020
rect 368584 4010 368612 330482
rect 368676 6458 368704 335326
rect 369228 316034 369256 338014
rect 369596 330546 369624 338014
rect 369584 330540 369636 330546
rect 369584 330482 369636 330488
rect 369860 323196 369912 323202
rect 369860 323138 369912 323144
rect 368768 316006 369256 316034
rect 368768 312594 368796 316006
rect 368756 312588 368808 312594
rect 368756 312530 368808 312536
rect 368756 18624 368808 18630
rect 368756 18566 368808 18572
rect 368768 16574 368796 18566
rect 368768 16546 369440 16574
rect 368664 6452 368716 6458
rect 368664 6394 368716 6400
rect 368572 4004 368624 4010
rect 368572 3946 368624 3952
rect 369412 480 369440 16546
rect 369872 3942 369900 323138
rect 369964 6390 369992 338014
rect 370332 318170 370360 338014
rect 370504 336320 370556 336326
rect 370504 336262 370556 336268
rect 370320 318164 370372 318170
rect 370320 318106 370372 318112
rect 370516 18630 370544 336262
rect 370700 323202 370728 338014
rect 371298 337770 371326 338028
rect 371528 338014 371680 338042
rect 371804 338014 372048 338042
rect 372172 338014 372416 338042
rect 372724 338014 372784 338042
rect 373092 338014 373152 338042
rect 373276 338014 373520 338042
rect 373644 338014 373888 338042
rect 374104 338014 374256 338042
rect 374380 338014 374624 338042
rect 374748 338014 374992 338042
rect 375300 338014 375360 338042
rect 375576 338014 375728 338042
rect 375852 338014 376096 338042
rect 376220 338014 376464 338042
rect 376832 338014 376984 338042
rect 371298 337742 371372 337770
rect 371240 326460 371292 326466
rect 371240 326402 371292 326408
rect 370688 323196 370740 323202
rect 370688 323138 370740 323144
rect 370504 18624 370556 18630
rect 370504 18566 370556 18572
rect 370596 9036 370648 9042
rect 370596 8978 370648 8984
rect 369952 6384 370004 6390
rect 369952 6326 370004 6332
rect 369860 3936 369912 3942
rect 369860 3878 369912 3884
rect 370608 480 370636 8978
rect 371252 3874 371280 326402
rect 371344 6322 371372 337742
rect 371424 325780 371476 325786
rect 371424 325722 371476 325728
rect 371332 6316 371384 6322
rect 371332 6258 371384 6264
rect 371436 6254 371464 325722
rect 371528 305726 371556 338014
rect 371804 326466 371832 338014
rect 371792 326460 371844 326466
rect 371792 326402 371844 326408
rect 372172 325786 372200 338014
rect 372620 326460 372672 326466
rect 372620 326402 372672 326408
rect 372160 325780 372212 325786
rect 372160 325722 372212 325728
rect 371516 305720 371568 305726
rect 371516 305662 371568 305668
rect 372632 10810 372660 326402
rect 372724 10878 372752 338014
rect 373092 336326 373120 338014
rect 373080 336320 373132 336326
rect 373080 336262 373132 336268
rect 373276 335354 373304 338014
rect 373356 336524 373408 336530
rect 373356 336466 373408 336472
rect 373184 335326 373304 335354
rect 373184 316034 373212 335326
rect 373368 316034 373396 336466
rect 373644 326466 373672 338014
rect 374000 336116 374052 336122
rect 374000 336058 374052 336064
rect 373632 326460 373684 326466
rect 373632 326402 373684 326408
rect 372816 316006 373212 316034
rect 373276 316006 373396 316034
rect 372816 279478 372844 316006
rect 372804 279472 372856 279478
rect 372804 279414 372856 279420
rect 372804 25560 372856 25566
rect 372804 25502 372856 25508
rect 372816 16574 372844 25502
rect 372816 16546 372936 16574
rect 372712 10872 372764 10878
rect 372712 10814 372764 10820
rect 372620 10804 372672 10810
rect 372620 10746 372672 10752
rect 371516 10328 371568 10334
rect 371516 10270 371568 10276
rect 371424 6248 371476 6254
rect 371424 6190 371476 6196
rect 371240 3868 371292 3874
rect 371240 3810 371292 3816
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371528 354 371556 10270
rect 372908 480 372936 16546
rect 373276 11762 373304 316006
rect 373264 11756 373316 11762
rect 373264 11698 373316 11704
rect 374012 3534 374040 336058
rect 374104 6914 374132 338014
rect 374184 326460 374236 326466
rect 374184 326402 374236 326408
rect 374196 10742 374224 326402
rect 374380 316034 374408 338014
rect 374748 326466 374776 338014
rect 375300 336258 375328 338014
rect 375288 336252 375340 336258
rect 375288 336194 375340 336200
rect 375576 326534 375604 338014
rect 375852 335354 375880 338014
rect 375668 335326 375880 335354
rect 375564 326528 375616 326534
rect 375564 326470 375616 326476
rect 374736 326460 374788 326466
rect 374736 326402 374788 326408
rect 375380 326460 375432 326466
rect 375380 326402 375432 326408
rect 374288 316006 374408 316034
rect 374288 278050 374316 316006
rect 374276 278044 374328 278050
rect 374276 277986 374328 277992
rect 374276 11824 374328 11830
rect 374276 11766 374328 11772
rect 374184 10736 374236 10742
rect 374184 10678 374236 10684
rect 374104 6886 374224 6914
rect 374196 3806 374224 6886
rect 374184 3800 374236 3806
rect 374184 3742 374236 3748
rect 374000 3528 374052 3534
rect 374288 3482 374316 11766
rect 375392 3738 375420 326402
rect 375668 321722 375696 335326
rect 375748 326528 375800 326534
rect 375748 326470 375800 326476
rect 375484 321694 375696 321722
rect 375484 10674 375512 321694
rect 375760 318794 375788 326470
rect 376220 326466 376248 338014
rect 376760 336728 376812 336734
rect 376760 336670 376812 336676
rect 376208 326460 376260 326466
rect 376208 326402 376260 326408
rect 375576 318766 375788 318794
rect 375576 276690 375604 318766
rect 375564 276684 375616 276690
rect 375564 276626 375616 276632
rect 375564 26920 375616 26926
rect 375564 26862 375616 26868
rect 375576 16574 375604 26862
rect 375576 16546 376064 16574
rect 375472 10668 375524 10674
rect 375472 10610 375524 10616
rect 375380 3732 375432 3738
rect 375380 3674 375432 3680
rect 374000 3470 374052 3476
rect 374104 3454 374316 3482
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 374104 480 374132 3454
rect 375300 480 375328 3470
rect 371670 354 371782 480
rect 371528 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 376772 10606 376800 336670
rect 376852 326460 376904 326466
rect 376852 326402 376904 326408
rect 376864 273970 376892 326402
rect 376956 275330 376984 338014
rect 377048 338014 377200 338042
rect 377508 338014 377568 338042
rect 377692 338014 377936 338042
rect 377048 336734 377076 338014
rect 377036 336728 377088 336734
rect 377036 336670 377088 336676
rect 377508 336190 377536 338014
rect 377496 336184 377548 336190
rect 377496 336126 377548 336132
rect 377404 336048 377456 336054
rect 377404 335990 377456 335996
rect 376944 275324 376996 275330
rect 376944 275266 376996 275272
rect 376852 273964 376904 273970
rect 376852 273906 376904 273912
rect 377312 13116 377364 13122
rect 377312 13058 377364 13064
rect 376760 10600 376812 10606
rect 376760 10542 376812 10548
rect 377324 3482 377352 13058
rect 377416 8294 377444 335990
rect 377692 326466 377720 338014
rect 378290 337770 378318 338028
rect 378428 338014 378672 338042
rect 378796 338014 379040 338042
rect 379164 338014 379316 338042
rect 379684 338014 379928 338042
rect 378290 337742 378364 337770
rect 378336 326738 378364 337742
rect 378324 326732 378376 326738
rect 378324 326674 378376 326680
rect 378428 326618 378456 338014
rect 378152 326590 378456 326618
rect 377680 326460 377732 326466
rect 377680 326402 377732 326408
rect 377404 8288 377456 8294
rect 377404 8230 377456 8236
rect 378152 3670 378180 326590
rect 378324 326528 378376 326534
rect 378324 326470 378376 326476
rect 378232 326460 378284 326466
rect 378232 326402 378284 326408
rect 378244 10470 378272 326402
rect 378336 10538 378364 326470
rect 378796 316034 378824 338014
rect 379164 326466 379192 338014
rect 379900 336122 379928 338014
rect 379992 338014 380052 338042
rect 380176 338014 380420 338042
rect 380544 338014 380788 338042
rect 381096 338014 381156 338042
rect 381280 338014 381524 338042
rect 381832 338014 381892 338042
rect 382016 338014 382260 338042
rect 382384 338014 382628 338042
rect 382752 338014 382996 338042
rect 383364 338014 383608 338042
rect 383732 338014 383884 338042
rect 379888 336116 379940 336122
rect 379888 336058 379940 336064
rect 379992 335442 380020 338014
rect 379980 335436 380032 335442
rect 379980 335378 380032 335384
rect 379152 326460 379204 326466
rect 379152 326402 379204 326408
rect 379520 326460 379572 326466
rect 379520 326402 379572 326408
rect 378428 316006 378824 316034
rect 378428 286346 378456 316006
rect 378416 286340 378468 286346
rect 378416 286282 378468 286288
rect 378324 10532 378376 10538
rect 378324 10474 378376 10480
rect 378232 10464 378284 10470
rect 378232 10406 378284 10412
rect 378876 8288 378928 8294
rect 378876 8230 378928 8236
rect 378140 3664 378192 3670
rect 378140 3606 378192 3612
rect 377324 3454 377720 3482
rect 377692 480 377720 3454
rect 378888 480 378916 8230
rect 379532 3534 379560 326402
rect 380176 316034 380204 338014
rect 380544 326466 380572 338014
rect 381096 326466 381124 338014
rect 381280 335354 381308 338014
rect 381832 336054 381860 338014
rect 381820 336048 381872 336054
rect 381820 335990 381872 335996
rect 381544 335436 381596 335442
rect 381544 335378 381596 335384
rect 381188 335326 381308 335354
rect 380532 326460 380584 326466
rect 380532 326402 380584 326408
rect 381084 326460 381136 326466
rect 381084 326402 381136 326408
rect 380900 322788 380952 322794
rect 380900 322730 380952 322736
rect 379624 316006 380204 316034
rect 379624 304298 379652 316006
rect 379612 304292 379664 304298
rect 379612 304234 379664 304240
rect 380912 7614 380940 322730
rect 381188 321858 381216 335326
rect 381268 326460 381320 326466
rect 381268 326402 381320 326408
rect 381004 321830 381216 321858
rect 381004 10402 381032 321830
rect 381280 318794 381308 326402
rect 381096 318766 381308 318794
rect 381096 284986 381124 318766
rect 381084 284980 381136 284986
rect 381084 284922 381136 284928
rect 381556 271182 381584 335378
rect 382016 322794 382044 338014
rect 382280 326460 382332 326466
rect 382280 326402 382332 326408
rect 382004 322788 382056 322794
rect 382004 322730 382056 322736
rect 381544 271176 381596 271182
rect 381544 271118 381596 271124
rect 381176 14476 381228 14482
rect 381176 14418 381228 14424
rect 380992 10396 381044 10402
rect 380992 10338 381044 10344
rect 379980 7608 380032 7614
rect 379980 7550 380032 7556
rect 380900 7608 380952 7614
rect 380900 7550 380952 7556
rect 379520 3528 379572 3534
rect 379520 3470 379572 3476
rect 379992 480 380020 7550
rect 381188 480 381216 14418
rect 382292 3505 382320 326402
rect 382384 10334 382412 338014
rect 382752 326466 382780 338014
rect 383014 336832 383070 336841
rect 383014 336767 383070 336776
rect 382924 336456 382976 336462
rect 382924 336398 382976 336404
rect 382740 326460 382792 326466
rect 382740 326402 382792 326408
rect 382464 21412 382516 21418
rect 382464 21354 382516 21360
rect 382372 10328 382424 10334
rect 382372 10270 382424 10276
rect 382476 6914 382504 21354
rect 382384 6886 382504 6914
rect 382278 3496 382334 3505
rect 382278 3431 382334 3440
rect 382384 480 382412 6886
rect 382936 4554 382964 336398
rect 383028 306338 383056 336767
rect 383580 334694 383608 338014
rect 383568 334688 383620 334694
rect 383568 334630 383620 334636
rect 383856 331226 383884 338014
rect 383948 338014 384100 338042
rect 383844 331220 383896 331226
rect 383844 331162 383896 331168
rect 383948 326754 383976 338014
rect 384454 337770 384482 338028
rect 384592 338014 384836 338042
rect 385144 338014 385204 338042
rect 385328 338014 385572 338042
rect 385696 338014 385940 338042
rect 386064 338014 386308 338042
rect 384454 337742 384528 337770
rect 384500 333334 384528 337742
rect 384488 333328 384540 333334
rect 384488 333270 384540 333276
rect 384028 331220 384080 331226
rect 384028 331162 384080 331168
rect 383672 326726 383976 326754
rect 383016 306332 383068 306338
rect 383016 306274 383068 306280
rect 383672 14482 383700 326726
rect 383752 326460 383804 326466
rect 383752 326402 383804 326408
rect 383764 268394 383792 326402
rect 384040 316034 384068 331162
rect 384592 326466 384620 338014
rect 384580 326460 384632 326466
rect 384580 326402 384632 326408
rect 385040 326324 385092 326330
rect 385040 326266 385092 326272
rect 383856 316006 384068 316034
rect 383856 269822 383884 316006
rect 383844 269816 383896 269822
rect 383844 269758 383896 269764
rect 383752 268388 383804 268394
rect 383752 268330 383804 268336
rect 385052 25566 385080 326266
rect 385144 247722 385172 338014
rect 385224 326460 385276 326466
rect 385224 326402 385276 326408
rect 385236 267034 385264 326402
rect 385328 320958 385356 338014
rect 385696 326466 385724 338014
rect 385684 326460 385736 326466
rect 385684 326402 385736 326408
rect 386064 326330 386092 338014
rect 386662 337770 386690 338028
rect 386800 338014 387044 338042
rect 387168 338014 387412 338042
rect 387536 338014 387780 338042
rect 387996 338014 388148 338042
rect 388272 338014 388516 338042
rect 388640 338014 388884 338042
rect 389192 338014 389252 338042
rect 389376 338014 389620 338042
rect 386662 337742 386736 337770
rect 386420 336728 386472 336734
rect 386420 336670 386472 336676
rect 386052 326324 386104 326330
rect 386052 326266 386104 326272
rect 385316 320952 385368 320958
rect 385316 320894 385368 320900
rect 385224 267028 385276 267034
rect 385224 266970 385276 266976
rect 386432 265674 386460 336670
rect 386512 326460 386564 326466
rect 386512 326402 386564 326408
rect 386420 265668 386472 265674
rect 386420 265610 386472 265616
rect 385132 247716 385184 247722
rect 385132 247658 385184 247664
rect 386524 246430 386552 326402
rect 386604 326324 386656 326330
rect 386604 326266 386656 326272
rect 386616 318102 386644 326266
rect 386708 319462 386736 337742
rect 386800 336734 386828 338014
rect 386788 336728 386840 336734
rect 386788 336670 386840 336676
rect 387064 336388 387116 336394
rect 387064 336330 387116 336336
rect 386696 319456 386748 319462
rect 386696 319398 386748 319404
rect 386604 318096 386656 318102
rect 386604 318038 386656 318044
rect 386512 246424 386564 246430
rect 386512 246366 386564 246372
rect 386420 246356 386472 246362
rect 386420 246298 386472 246304
rect 385132 47592 385184 47598
rect 385132 47534 385184 47540
rect 385040 25560 385092 25566
rect 385040 25502 385092 25508
rect 385144 16574 385172 47534
rect 386432 16574 386460 246298
rect 385144 16546 386000 16574
rect 386432 16546 386736 16574
rect 383660 14476 383712 14482
rect 383660 14418 383712 14424
rect 383568 8968 383620 8974
rect 383568 8910 383620 8916
rect 382924 4548 382976 4554
rect 382924 4490 382976 4496
rect 383580 480 383608 8910
rect 384764 4548 384816 4554
rect 384764 4490 384816 4496
rect 384776 480 384804 4490
rect 385972 480 386000 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387076 8974 387104 336330
rect 387168 326466 387196 338014
rect 387156 326460 387208 326466
rect 387156 326402 387208 326408
rect 387536 326330 387564 338014
rect 387800 326460 387852 326466
rect 387800 326402 387852 326408
rect 387524 326324 387576 326330
rect 387524 326266 387576 326272
rect 387812 316742 387840 326402
rect 387892 322176 387944 322182
rect 387892 322118 387944 322124
rect 387800 316736 387852 316742
rect 387800 316678 387852 316684
rect 387800 286408 387852 286414
rect 387800 286350 387852 286356
rect 387064 8968 387116 8974
rect 387064 8910 387116 8916
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 286350
rect 387904 243574 387932 322118
rect 387996 264246 388024 338014
rect 388272 322182 388300 338014
rect 388640 326466 388668 338014
rect 388628 326460 388680 326466
rect 388628 326402 388680 326408
rect 388260 322176 388312 322182
rect 388260 322118 388312 322124
rect 387984 264240 388036 264246
rect 387984 264182 388036 264188
rect 389192 262886 389220 338014
rect 389376 335354 389404 338014
rect 389974 337770 390002 338028
rect 390112 338014 390356 338042
rect 390664 338014 390724 338042
rect 390848 338014 391092 338042
rect 391216 338014 391368 338042
rect 391492 338014 391736 338042
rect 389974 337742 390048 337770
rect 389284 335326 389404 335354
rect 389180 262880 389232 262886
rect 389180 262822 389232 262828
rect 389180 261520 389232 261526
rect 389180 261462 389232 261468
rect 387892 243568 387944 243574
rect 387892 243510 387944 243516
rect 389192 16574 389220 261462
rect 389284 242214 389312 335326
rect 390020 331974 390048 337742
rect 390008 331968 390060 331974
rect 390008 331910 390060 331916
rect 390112 316034 390140 338014
rect 390560 330472 390612 330478
rect 390560 330414 390612 330420
rect 389376 316006 390140 316034
rect 389376 261526 389404 316006
rect 389364 261520 389416 261526
rect 389364 261462 389416 261468
rect 389272 242208 389324 242214
rect 389272 242150 389324 242156
rect 390572 26926 390600 330414
rect 390664 240786 390692 338014
rect 390744 330540 390796 330546
rect 390744 330482 390796 330488
rect 390756 283626 390784 330482
rect 390848 305658 390876 338014
rect 391216 330546 391244 338014
rect 391204 330540 391256 330546
rect 391204 330482 391256 330488
rect 391492 330478 391520 338014
rect 392090 337770 392118 338028
rect 392228 338014 392472 338042
rect 392596 338014 392840 338042
rect 392964 338014 393208 338042
rect 393516 338014 393576 338042
rect 393700 338014 393944 338042
rect 394068 338014 394312 338042
rect 394436 338014 394680 338042
rect 394804 338014 395048 338042
rect 395172 338014 395416 338042
rect 395540 338014 395784 338042
rect 396152 338014 396304 338042
rect 392090 337742 392164 337770
rect 392032 330540 392084 330546
rect 392032 330482 392084 330488
rect 391480 330472 391532 330478
rect 391480 330414 391532 330420
rect 391940 330472 391992 330478
rect 391940 330414 391992 330420
rect 391952 313954 391980 330414
rect 391940 313948 391992 313954
rect 391940 313890 391992 313896
rect 390836 305652 390888 305658
rect 390836 305594 390888 305600
rect 390744 283620 390796 283626
rect 390744 283562 390796 283568
rect 391940 260160 391992 260166
rect 391940 260102 391992 260108
rect 390652 240780 390704 240786
rect 390652 240722 390704 240728
rect 390744 29640 390796 29646
rect 390744 29582 390796 29588
rect 390560 26920 390612 26926
rect 390560 26862 390612 26868
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390756 6914 390784 29582
rect 391952 16574 391980 260102
rect 392044 239426 392072 330482
rect 392136 329118 392164 337742
rect 392124 329112 392176 329118
rect 392124 329054 392176 329060
rect 392228 316034 392256 338014
rect 392596 330546 392624 338014
rect 392584 330540 392636 330546
rect 392584 330482 392636 330488
rect 392964 330478 392992 338014
rect 393412 330540 393464 330546
rect 393412 330482 393464 330488
rect 392952 330472 393004 330478
rect 392952 330414 393004 330420
rect 393320 327616 393372 327622
rect 393320 327558 393372 327564
rect 392136 316006 392256 316034
rect 392136 260166 392164 316006
rect 392124 260160 392176 260166
rect 392124 260102 392176 260108
rect 392032 239420 392084 239426
rect 392032 239362 392084 239368
rect 393332 28286 393360 327558
rect 393424 257378 393452 330482
rect 393516 301510 393544 338014
rect 393700 327622 393728 338014
rect 394068 327758 394096 338014
rect 394436 330546 394464 338014
rect 394424 330540 394476 330546
rect 394424 330482 394476 330488
rect 394700 329928 394752 329934
rect 394700 329870 394752 329876
rect 394056 327752 394108 327758
rect 394056 327694 394108 327700
rect 393688 327616 393740 327622
rect 393688 327558 393740 327564
rect 394712 315314 394740 329870
rect 394700 315308 394752 315314
rect 394700 315250 394752 315256
rect 393504 301504 393556 301510
rect 393504 301446 393556 301452
rect 394700 285048 394752 285054
rect 394700 284990 394752 284996
rect 393412 257372 393464 257378
rect 393412 257314 393464 257320
rect 393412 28416 393464 28422
rect 393412 28358 393464 28364
rect 393320 28280 393372 28286
rect 393320 28222 393372 28228
rect 393424 16574 393452 28358
rect 394712 16574 394740 284990
rect 394804 238066 394832 338014
rect 395172 329934 395200 338014
rect 395160 329928 395212 329934
rect 395160 329870 395212 329876
rect 395540 316034 395568 338014
rect 396080 330540 396132 330546
rect 396080 330482 396132 330488
rect 394896 316006 395568 316034
rect 394896 282198 394924 316006
rect 394884 282192 394936 282198
rect 394884 282134 394936 282140
rect 394792 238060 394844 238066
rect 394792 238002 394844 238008
rect 396092 21418 396120 330482
rect 396172 330472 396224 330478
rect 396172 330414 396224 330420
rect 396184 235278 396212 330414
rect 396276 236706 396304 338014
rect 396460 338014 396520 338042
rect 396644 338014 396888 338042
rect 397012 338014 397256 338042
rect 397624 338014 397776 338042
rect 396460 336394 396488 338014
rect 396448 336388 396500 336394
rect 396448 336330 396500 336336
rect 396644 330546 396672 338014
rect 396632 330540 396684 330546
rect 396632 330482 396684 330488
rect 397012 330478 397040 338014
rect 397552 336728 397604 336734
rect 397552 336670 397604 336676
rect 397000 330472 397052 330478
rect 397000 330414 397052 330420
rect 397460 330472 397512 330478
rect 397460 330414 397512 330420
rect 396264 236700 396316 236706
rect 396264 236642 396316 236648
rect 396172 235272 396224 235278
rect 396172 235214 396224 235220
rect 397472 233918 397500 330414
rect 397564 300150 397592 336670
rect 397644 330540 397696 330546
rect 397644 330482 397696 330488
rect 397656 322250 397684 330482
rect 397748 323610 397776 338014
rect 397840 338014 397992 338042
rect 398116 338014 398360 338042
rect 398484 338014 398728 338042
rect 398944 338014 399096 338042
rect 399220 338014 399464 338042
rect 399772 338014 399832 338042
rect 399956 338014 400200 338042
rect 400324 338014 400568 338042
rect 400692 338014 400936 338042
rect 401060 338014 401304 338042
rect 401672 338014 401824 338042
rect 397840 336734 397868 338014
rect 397828 336728 397880 336734
rect 397828 336670 397880 336676
rect 398116 330478 398144 338014
rect 398484 330546 398512 338014
rect 398472 330540 398524 330546
rect 398472 330482 398524 330488
rect 398104 330472 398156 330478
rect 398104 330414 398156 330420
rect 398944 326466 398972 338014
rect 399220 331214 399248 338014
rect 399772 336598 399800 338014
rect 399760 336592 399812 336598
rect 399760 336534 399812 336540
rect 399036 331186 399248 331214
rect 398932 326460 398984 326466
rect 398932 326402 398984 326408
rect 397736 323604 397788 323610
rect 397736 323546 397788 323552
rect 397644 322244 397696 322250
rect 397644 322186 397696 322192
rect 399036 321722 399064 331186
rect 399116 326460 399168 326466
rect 399116 326402 399168 326408
rect 398852 321694 399064 321722
rect 397552 300144 397604 300150
rect 397552 300086 397604 300092
rect 397460 233912 397512 233918
rect 397460 233854 397512 233860
rect 398852 42090 398880 321694
rect 399128 318794 399156 326402
rect 398944 318766 399156 318794
rect 398944 291854 398972 318766
rect 399956 316034 399984 338014
rect 400324 336682 400352 338014
rect 399036 316006 399984 316034
rect 400232 336654 400352 336682
rect 398932 291848 398984 291854
rect 398932 291790 398984 291796
rect 399036 256018 399064 316006
rect 398932 256012 398984 256018
rect 398932 255954 398984 255960
rect 399024 256012 399076 256018
rect 399024 255954 399076 255960
rect 398840 42084 398892 42090
rect 398840 42026 398892 42032
rect 397460 32428 397512 32434
rect 397460 32370 397512 32376
rect 396172 22772 396224 22778
rect 396172 22714 396224 22720
rect 396080 21412 396132 21418
rect 396080 21354 396132 21360
rect 391952 16546 392624 16574
rect 393424 16546 394280 16574
rect 394712 16546 395384 16574
rect 390664 6886 390784 6914
rect 390664 480 390692 6886
rect 391848 4820 391900 4826
rect 391848 4762 391900 4768
rect 391860 480 391888 4762
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396184 354 396212 22714
rect 397472 16574 397500 32370
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398840 8968 398892 8974
rect 398840 8910 398892 8916
rect 398852 3074 398880 8910
rect 398944 3194 398972 255954
rect 400232 32434 400260 336654
rect 400692 335354 400720 338014
rect 401060 336682 401088 338014
rect 400324 335326 400720 335354
rect 400784 336654 401088 336682
rect 401600 336728 401652 336734
rect 401600 336670 401652 336676
rect 400324 297430 400352 335326
rect 400784 316034 400812 336654
rect 400864 336592 400916 336598
rect 400864 336534 400916 336540
rect 400416 316006 400812 316034
rect 400312 297424 400364 297430
rect 400312 297366 400364 297372
rect 400416 254590 400444 316006
rect 400876 311166 400904 336534
rect 400864 311160 400916 311166
rect 400864 311102 400916 311108
rect 400312 254584 400364 254590
rect 400312 254526 400364 254532
rect 400404 254584 400456 254590
rect 400404 254526 400456 254532
rect 400220 32428 400272 32434
rect 400220 32370 400272 32376
rect 400324 16574 400352 254526
rect 400324 16546 400904 16574
rect 398932 3188 398984 3194
rect 398932 3130 398984 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396184 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 401612 4826 401640 336670
rect 401692 326460 401744 326466
rect 401692 326402 401744 326408
rect 401704 229770 401732 326402
rect 401796 231130 401824 338014
rect 401888 338014 402040 338042
rect 402348 338014 402408 338042
rect 402532 338014 402776 338042
rect 401888 336734 401916 338014
rect 401876 336728 401928 336734
rect 401876 336670 401928 336676
rect 402348 335374 402376 338014
rect 402336 335368 402388 335374
rect 402336 335310 402388 335316
rect 402532 326466 402560 338014
rect 403130 337770 403158 338028
rect 403268 338014 403420 338042
rect 403130 337742 403204 337770
rect 403176 334626 403204 337742
rect 403164 334620 403216 334626
rect 403164 334562 403216 334568
rect 403268 331214 403296 338014
rect 403774 337770 403802 338028
rect 403912 338014 404156 338042
rect 404464 338014 404524 338042
rect 404648 338014 404892 338042
rect 403774 337742 403848 337770
rect 403624 335368 403676 335374
rect 403624 335310 403676 335316
rect 402992 331186 403296 331214
rect 402520 326460 402572 326466
rect 402520 326402 402572 326408
rect 402992 290494 403020 331186
rect 403072 326460 403124 326466
rect 403072 326402 403124 326408
rect 403084 296002 403112 326402
rect 403072 295996 403124 296002
rect 403072 295938 403124 295944
rect 402980 290488 403032 290494
rect 402980 290430 403032 290436
rect 402980 272536 403032 272542
rect 402980 272478 403032 272484
rect 401784 231124 401836 231130
rect 401784 231066 401836 231072
rect 401692 229764 401744 229770
rect 401692 229706 401744 229712
rect 402992 16574 403020 272478
rect 403636 222902 403664 335310
rect 403820 331906 403848 337742
rect 403808 331900 403860 331906
rect 403808 331842 403860 331848
rect 403912 326466 403940 338014
rect 404464 326466 404492 338014
rect 404648 335354 404676 338014
rect 405246 337770 405274 338028
rect 405384 338014 405628 338042
rect 405844 338014 405996 338042
rect 406120 338014 406364 338042
rect 406488 338014 406732 338042
rect 406856 338014 407100 338042
rect 407316 338014 407468 338042
rect 407592 338014 407836 338042
rect 407960 338014 408204 338042
rect 408512 338014 408572 338042
rect 408696 338014 408940 338042
rect 409064 338014 409308 338042
rect 409432 338014 409676 338042
rect 405246 337742 405320 337770
rect 404556 335326 404676 335354
rect 403900 326460 403952 326466
rect 403900 326402 403952 326408
rect 404452 326460 404504 326466
rect 404452 326402 404504 326408
rect 404556 321722 404584 335326
rect 405292 330410 405320 337742
rect 405280 330404 405332 330410
rect 405280 330346 405332 330352
rect 404636 326460 404688 326466
rect 404636 326402 404688 326408
rect 404372 321694 404584 321722
rect 403624 222896 403676 222902
rect 403624 222838 403676 222844
rect 402992 16546 403664 16574
rect 402520 15904 402572 15910
rect 402520 15846 402572 15852
rect 401600 4820 401652 4826
rect 401600 4762 401652 4768
rect 402532 480 402560 15846
rect 403636 480 403664 16546
rect 404372 15910 404400 321694
rect 404648 318794 404676 326402
rect 404464 318766 404676 318794
rect 404464 253230 404492 318766
rect 405384 316034 405412 338014
rect 405740 326324 405792 326330
rect 405740 326266 405792 326272
rect 404556 316006 405412 316034
rect 404556 280838 404584 316006
rect 404544 280832 404596 280838
rect 404544 280774 404596 280780
rect 404452 253224 404504 253230
rect 404452 253166 404504 253172
rect 404452 31068 404504 31074
rect 404452 31010 404504 31016
rect 404360 15904 404412 15910
rect 404360 15846 404412 15852
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404464 354 404492 31010
rect 405752 17270 405780 326266
rect 405844 228410 405872 338014
rect 405924 326460 405976 326466
rect 405924 326402 405976 326408
rect 405936 289134 405964 326402
rect 406120 316034 406148 338014
rect 406488 326466 406516 338014
rect 406476 326460 406528 326466
rect 406476 326402 406528 326408
rect 406856 326330 406884 338014
rect 407120 326460 407172 326466
rect 407120 326402 407172 326408
rect 406844 326324 406896 326330
rect 406844 326266 406896 326272
rect 406028 316006 406148 316034
rect 406028 309806 406056 316006
rect 406016 309800 406068 309806
rect 406016 309742 406068 309748
rect 405924 289128 405976 289134
rect 405924 289070 405976 289076
rect 405832 228404 405884 228410
rect 405832 228346 405884 228352
rect 405832 17400 405884 17406
rect 405832 17342 405884 17348
rect 405740 17264 405792 17270
rect 405740 17206 405792 17212
rect 405844 16574 405872 17342
rect 405844 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 13122 407160 326402
rect 407212 324284 407264 324290
rect 407212 324226 407264 324232
rect 407224 227050 407252 324226
rect 407316 294642 407344 338014
rect 407592 326466 407620 338014
rect 407580 326460 407632 326466
rect 407580 326402 407632 326408
rect 407960 324290 407988 338014
rect 408512 333266 408540 338014
rect 408500 333260 408552 333266
rect 408500 333202 408552 333208
rect 408500 324556 408552 324562
rect 408500 324498 408552 324504
rect 407948 324284 408000 324290
rect 407948 324226 408000 324232
rect 407304 294636 407356 294642
rect 407304 294578 407356 294584
rect 407212 227044 407264 227050
rect 407212 226986 407264 226992
rect 408512 29646 408540 324498
rect 408592 323876 408644 323882
rect 408592 323818 408644 323824
rect 408604 308446 408632 323818
rect 408592 308440 408644 308446
rect 408592 308382 408644 308388
rect 408592 283688 408644 283694
rect 408592 283630 408644 283636
rect 408500 29640 408552 29646
rect 408500 29582 408552 29588
rect 407212 24132 407264 24138
rect 407212 24074 407264 24080
rect 407120 13116 407172 13122
rect 407120 13058 407172 13064
rect 407224 480 407252 24074
rect 408604 16574 408632 283630
rect 408696 251870 408724 338014
rect 409064 324562 409092 338014
rect 409052 324556 409104 324562
rect 409052 324498 409104 324504
rect 409432 323882 409460 338014
rect 410030 337770 410058 338028
rect 410260 338014 410412 338042
rect 410536 338014 410780 338042
rect 410904 338014 411148 338042
rect 411272 338014 411516 338042
rect 411824 338014 411884 338042
rect 412008 338014 412252 338042
rect 412376 338014 412620 338042
rect 412744 338014 412988 338042
rect 413112 338014 413356 338042
rect 413480 338014 413724 338042
rect 410030 337742 410104 337770
rect 410076 326534 410104 337742
rect 410064 326528 410116 326534
rect 410064 326470 410116 326476
rect 409880 326460 409932 326466
rect 409880 326402 409932 326408
rect 409420 323876 409472 323882
rect 409420 323818 409472 323824
rect 409892 307086 409920 326402
rect 410260 326346 410288 338014
rect 410340 326528 410392 326534
rect 410340 326470 410392 326476
rect 409984 326318 410288 326346
rect 409880 307080 409932 307086
rect 409880 307022 409932 307028
rect 408684 251864 408736 251870
rect 408684 251806 408736 251812
rect 409880 250504 409932 250510
rect 409880 250446 409932 250452
rect 409892 16574 409920 250446
rect 409984 225622 410012 326318
rect 410064 326256 410116 326262
rect 410064 326198 410116 326204
rect 410076 249082 410104 326198
rect 410352 321554 410380 326470
rect 410536 326466 410564 338014
rect 410524 326460 410576 326466
rect 410524 326402 410576 326408
rect 410904 326262 410932 338014
rect 410892 326256 410944 326262
rect 410892 326198 410944 326204
rect 410168 321526 410380 321554
rect 410168 250510 410196 321526
rect 410156 250504 410208 250510
rect 410156 250446 410208 250452
rect 410064 249076 410116 249082
rect 410064 249018 410116 249024
rect 409972 225616 410024 225622
rect 409972 225558 410024 225564
rect 411272 36582 411300 338014
rect 411824 335374 411852 338014
rect 411812 335368 411864 335374
rect 411812 335310 411864 335316
rect 411352 326460 411404 326466
rect 411352 326402 411404 326408
rect 411364 224262 411392 326402
rect 412008 316034 412036 338014
rect 412376 326466 412404 338014
rect 412744 334642 412772 338014
rect 412652 334614 412772 334642
rect 412364 326460 412416 326466
rect 412364 326402 412416 326408
rect 411456 316006 412036 316034
rect 411456 287706 411484 316006
rect 411444 287700 411496 287706
rect 411444 287642 411496 287648
rect 411352 224256 411404 224262
rect 411352 224198 411404 224204
rect 411260 36576 411312 36582
rect 411260 36518 411312 36524
rect 408604 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 3596 408460 3602
rect 408408 3538 408460 3544
rect 408420 480 408448 3538
rect 404790 354 404902 480
rect 404464 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 412652 6186 412680 334614
rect 413112 331214 413140 338014
rect 413480 335458 413508 338014
rect 414078 337770 414106 338028
rect 414216 338014 414460 338042
rect 414584 338014 414828 338042
rect 414078 337742 414152 337770
rect 412744 331186 413140 331214
rect 413204 335430 413508 335458
rect 412744 8974 412772 331186
rect 413204 320890 413232 335430
rect 413376 335368 413428 335374
rect 413376 335310 413428 335316
rect 413388 331214 413416 335310
rect 414020 334552 414072 334558
rect 414020 334494 414072 334500
rect 413296 331186 413416 331214
rect 413192 320884 413244 320890
rect 413192 320826 413244 320832
rect 413296 293282 413324 331186
rect 413284 293276 413336 293282
rect 413284 293218 413336 293224
rect 412824 18624 412876 18630
rect 412824 18566 412876 18572
rect 412732 8968 412784 8974
rect 412732 8910 412784 8916
rect 412640 6180 412692 6186
rect 412640 6122 412692 6128
rect 411904 3460 411956 3466
rect 411904 3402 411956 3408
rect 411916 480 411944 3402
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412836 354 412864 18566
rect 414032 3194 414060 334494
rect 414124 3602 414152 337742
rect 414216 334558 414244 338014
rect 414204 334552 414256 334558
rect 414204 334494 414256 334500
rect 414584 316034 414612 338014
rect 414216 316006 414612 316034
rect 414112 3596 414164 3602
rect 414112 3538 414164 3544
rect 414216 3369 414244 316006
rect 414952 20670 414980 457422
rect 416780 324964 416832 324970
rect 416780 324906 416832 324912
rect 415400 282260 415452 282266
rect 415400 282202 415452 282208
rect 414940 20664 414992 20670
rect 414940 20606 414992 20612
rect 414296 11756 414348 11762
rect 414296 11698 414348 11704
rect 414202 3360 414258 3369
rect 414202 3295 414258 3304
rect 414020 3188 414072 3194
rect 414020 3130 414072 3136
rect 414308 480 414336 11698
rect 415412 3466 415440 282202
rect 416792 16574 416820 324906
rect 417436 46918 417464 458322
rect 417528 431934 417556 461246
rect 422944 461236 422996 461242
rect 422944 461178 422996 461184
rect 420184 461168 420236 461174
rect 420184 461110 420236 461116
rect 418804 458448 418856 458454
rect 418804 458390 418856 458396
rect 417516 431928 417568 431934
rect 417516 431870 417568 431876
rect 418816 86970 418844 458390
rect 420196 353258 420224 461110
rect 421564 458516 421616 458522
rect 421564 458458 421616 458464
rect 420184 353252 420236 353258
rect 420184 353194 420236 353200
rect 420182 331800 420238 331809
rect 420182 331735 420238 331744
rect 419540 326392 419592 326398
rect 419540 326334 419592 326340
rect 418804 86964 418856 86970
rect 418804 86906 418856 86912
rect 417424 46912 417476 46918
rect 417424 46854 417476 46860
rect 419552 16574 419580 326334
rect 420196 126954 420224 331735
rect 420920 321020 420972 321026
rect 420920 320962 420972 320968
rect 420184 126948 420236 126954
rect 420184 126890 420236 126896
rect 416792 16546 417464 16574
rect 419552 16546 420224 16574
rect 415492 13184 415544 13190
rect 415492 13126 415544 13132
rect 415400 3460 415452 3466
rect 415400 3402 415452 3408
rect 415504 480 415532 13126
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 416780 3460 416832 3466
rect 416780 3402 416832 3408
rect 416700 480 416728 3402
rect 416792 3194 416820 3402
rect 416780 3188 416832 3194
rect 416780 3130 416832 3136
rect 413070 354 413182 480
rect 412836 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418988 3256 419040 3262
rect 418988 3198 419040 3204
rect 419000 480 419028 3198
rect 420196 480 420224 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 320962
rect 421576 167006 421604 458458
rect 422956 405686 422984 461178
rect 462332 460766 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 460760 462372 460766
rect 462320 460702 462372 460708
rect 477512 460698 477540 702406
rect 494072 461650 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 461644 494112 461650
rect 494060 461586 494112 461592
rect 477500 460692 477552 460698
rect 477500 460634 477552 460640
rect 527192 460562 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 460556 527232 460562
rect 527180 460498 527232 460504
rect 542372 460494 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 542360 460488 542412 460494
rect 542360 460430 542412 460436
rect 424324 458788 424376 458794
rect 424324 458730 424376 458736
rect 422944 405680 422996 405686
rect 422944 405622 422996 405628
rect 424336 379506 424364 458730
rect 425704 458720 425756 458726
rect 425704 458662 425756 458668
rect 424324 379500 424376 379506
rect 424324 379442 424376 379448
rect 425716 365702 425744 458662
rect 580264 458312 580316 458318
rect 580264 458254 580316 458260
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 427084 456884 427136 456890
rect 427084 456826 427136 456832
rect 427096 419490 427124 456826
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 427084 419484 427136 419490
rect 427084 419426 427136 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 425704 365696 425756 365702
rect 425704 365638 425756 365644
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 422944 336388 422996 336394
rect 422944 336330 422996 336336
rect 421564 167000 421616 167006
rect 421564 166942 421616 166948
rect 422956 11762 422984 336330
rect 447140 336320 447192 336326
rect 447140 336262 447192 336268
rect 423680 330608 423732 330614
rect 423680 330550 423732 330556
rect 423034 329080 423090 329089
rect 423034 329015 423090 329024
rect 423048 245614 423076 329015
rect 423036 245608 423088 245614
rect 423036 245550 423088 245556
rect 422944 11756 422996 11762
rect 422944 11698 422996 11704
rect 422576 3324 422628 3330
rect 422576 3266 422628 3272
rect 422588 480 422616 3266
rect 423692 1018 423720 330550
rect 424322 327720 424378 327729
rect 424322 327655 424378 327664
rect 424336 299470 424364 327655
rect 425702 323640 425758 323649
rect 425702 323575 425758 323584
rect 424324 299464 424376 299470
rect 424324 299406 424376 299412
rect 423772 298784 423824 298790
rect 423772 298726 423824 298732
rect 423680 1012 423732 1018
rect 423680 954 423732 960
rect 423784 480 423812 298726
rect 424322 291816 424378 291825
rect 424322 291751 424378 291760
rect 424336 139398 424364 291751
rect 424324 139392 424376 139398
rect 424324 139334 424376 139340
rect 425716 73166 425744 323575
rect 438122 322144 438178 322153
rect 438122 322079 438178 322088
rect 427820 319524 427872 319530
rect 427820 319466 427872 319472
rect 427082 309768 427138 309777
rect 427082 309703 427138 309712
rect 426440 280900 426492 280906
rect 426440 280842 426492 280848
rect 425704 73160 425756 73166
rect 425704 73102 425756 73108
rect 426452 16574 426480 280842
rect 427096 153202 427124 309703
rect 427084 153196 427136 153202
rect 427084 153138 427136 153144
rect 427832 16574 427860 319466
rect 434720 312588 434772 312594
rect 434720 312530 434772 312536
rect 428462 308408 428518 308417
rect 428462 308343 428518 308352
rect 428476 193186 428504 308343
rect 429842 307048 429898 307057
rect 429842 306983 429898 306992
rect 429856 233238 429884 306983
rect 431222 301472 431278 301481
rect 431222 301407 431278 301416
rect 429844 233232 429896 233238
rect 429844 233174 429896 233180
rect 428464 193180 428516 193186
rect 428464 193122 428516 193128
rect 431236 60722 431264 301407
rect 432602 300112 432658 300121
rect 432602 300047 432658 300056
rect 432052 258732 432104 258738
rect 432052 258674 432104 258680
rect 431224 60716 431276 60722
rect 431224 60658 431276 60664
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 426164 3392 426216 3398
rect 426164 3334 426216 3340
rect 424968 1012 425020 1018
rect 424968 954 425020 960
rect 424980 480 425008 954
rect 426176 480 426204 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 430856 6520 430908 6526
rect 430856 6462 430908 6468
rect 429660 4140 429712 4146
rect 429660 4082 429712 4088
rect 429672 480 429700 4082
rect 430868 480 430896 6462
rect 432064 480 432092 258674
rect 432616 100706 432644 300047
rect 432604 100700 432656 100706
rect 432604 100642 432656 100648
rect 434732 16574 434760 312530
rect 435362 290456 435418 290465
rect 435362 290391 435418 290400
rect 435376 179382 435404 290391
rect 436742 289096 436798 289105
rect 436742 289031 436798 289040
rect 436756 219434 436784 289031
rect 436744 219428 436796 219434
rect 436744 219370 436796 219376
rect 435364 179376 435416 179382
rect 435364 179318 435416 179324
rect 438136 113150 438164 322079
rect 438860 318164 438912 318170
rect 438860 318106 438912 318112
rect 438124 113144 438176 113150
rect 438124 113086 438176 113092
rect 438872 16574 438900 318106
rect 441620 305720 441672 305726
rect 441620 305662 441672 305668
rect 441632 16574 441660 305662
rect 445022 287736 445078 287745
rect 445022 287671 445078 287680
rect 445036 259418 445064 287671
rect 445024 259412 445076 259418
rect 445024 259354 445076 259360
rect 447152 16574 447180 336262
rect 454040 336252 454092 336258
rect 454040 336194 454092 336200
rect 448520 279472 448572 279478
rect 448520 279414 448572 279420
rect 434732 16546 435128 16574
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 447152 16546 447456 16574
rect 434444 6452 434496 6458
rect 434444 6394 434496 6400
rect 433248 4072 433300 4078
rect 433248 4014 433300 4020
rect 433260 480 433288 4014
rect 434456 480 434484 6394
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 437940 6384 437992 6390
rect 437940 6326 437992 6332
rect 436744 4004 436796 4010
rect 436744 3946 436796 3952
rect 436756 480 436784 3946
rect 437952 480 437980 6326
rect 439148 480 439176 16546
rect 441528 6316 441580 6322
rect 441528 6258 441580 6264
rect 440332 3936 440384 3942
rect 440332 3878 440384 3884
rect 440344 480 440372 3878
rect 441540 480 441568 6258
rect 442644 480 442672 16546
rect 445760 10872 445812 10878
rect 445760 10814 445812 10820
rect 445024 6248 445076 6254
rect 445024 6190 445076 6196
rect 443828 3868 443880 3874
rect 443828 3810 443880 3816
rect 443840 480 443868 3810
rect 445036 480 445064 6190
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 10814
rect 447428 480 447456 16546
rect 448532 3210 448560 279414
rect 451280 278044 451332 278050
rect 451280 277986 451332 277992
rect 451292 16574 451320 277986
rect 451292 16546 451688 16574
rect 448612 10804 448664 10810
rect 448612 10746 448664 10752
rect 448624 3398 448652 10746
rect 450912 3800 450964 3806
rect 450912 3742 450964 3748
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 3742
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453304 10736 453356 10742
rect 453304 10678 453356 10684
rect 453316 480 453344 10678
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 336194
rect 460940 336184 460992 336190
rect 460940 336126 460992 336132
rect 460202 304192 460258 304201
rect 460202 304127 460258 304136
rect 455420 276684 455472 276690
rect 455420 276626 455472 276632
rect 455432 16574 455460 276626
rect 458180 275324 458232 275330
rect 458180 275266 458232 275272
rect 458192 16574 458220 275266
rect 460216 273222 460244 304127
rect 460204 273216 460256 273222
rect 460204 273158 460256 273164
rect 460952 16574 460980 336126
rect 467840 336116 467892 336122
rect 467840 336058 467892 336064
rect 465172 286340 465224 286346
rect 465172 286282 465224 286288
rect 462320 273964 462372 273970
rect 462320 273906 462372 273912
rect 455432 16546 455736 16574
rect 458192 16546 459232 16574
rect 460952 16546 461624 16574
rect 455708 480 455736 16546
rect 456892 10668 456944 10674
rect 456892 10610 456944 10616
rect 456904 480 456932 10610
rect 458088 3732 458140 3738
rect 458088 3674 458140 3680
rect 458100 480 458128 3674
rect 459204 480 459232 16546
rect 459928 10600 459980 10606
rect 459928 10542 459980 10548
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 10542
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 273906
rect 465184 16574 465212 286282
rect 467852 16574 467880 336058
rect 474740 336048 474792 336054
rect 474740 335990 474792 335996
rect 470600 304292 470652 304298
rect 470600 304234 470652 304240
rect 469220 271176 469272 271182
rect 469220 271118 469272 271124
rect 469232 16574 469260 271118
rect 465184 16546 465856 16574
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 463976 10532 464028 10538
rect 463976 10474 464028 10480
rect 463988 480 464016 10474
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 465184 480 465212 3606
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467472 10464 467524 10470
rect 467472 10406 467524 10412
rect 467484 480 467512 10406
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 304234
rect 473360 284980 473412 284986
rect 473360 284922 473412 284928
rect 473372 16574 473400 284922
rect 474752 16574 474780 335990
rect 480260 334688 480312 334694
rect 480260 334630 480312 334636
rect 479522 330440 479578 330449
rect 479522 330375 479578 330384
rect 479536 206990 479564 330375
rect 479524 206984 479576 206990
rect 479524 206926 479576 206932
rect 480272 16574 480300 334630
rect 543740 334620 543792 334626
rect 543740 334562 543792 334568
rect 483020 333328 483072 333334
rect 483020 333270 483072 333276
rect 481640 269816 481692 269822
rect 481640 269758 481692 269764
rect 481652 16574 481680 269758
rect 483032 16574 483060 333270
rect 500960 331968 501012 331974
rect 500960 331910 501012 331916
rect 487160 320952 487212 320958
rect 487160 320894 487212 320900
rect 484400 268388 484452 268394
rect 484400 268330 484452 268336
rect 484412 16574 484440 268330
rect 485780 247716 485832 247722
rect 485780 247658 485832 247664
rect 485792 16574 485820 247658
rect 473372 16546 473492 16574
rect 474752 16546 475792 16574
rect 480272 16546 480576 16574
rect 481652 16546 481772 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 472256 3528 472308 3534
rect 472256 3470 472308 3476
rect 472268 480 472296 3470
rect 473464 480 473492 16546
rect 474096 10396 474148 10402
rect 474096 10338 474148 10344
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 10338
rect 475764 480 475792 16546
rect 478144 10328 478196 10334
rect 478144 10270 478196 10276
rect 476948 7608 477000 7614
rect 476948 7550 477000 7556
rect 476960 480 476988 7550
rect 478156 480 478184 10270
rect 479338 3496 479394 3505
rect 479338 3431 479394 3440
rect 479352 480 479380 3431
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 482376 14476 482428 14482
rect 482376 14418 482428 14424
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 14418
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 320894
rect 489920 319456 489972 319462
rect 489920 319398 489972 319404
rect 488540 267028 488592 267034
rect 488540 266970 488592 266976
rect 488552 16574 488580 266970
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3534 489960 319398
rect 494060 318096 494112 318102
rect 494060 318038 494112 318044
rect 491300 265668 491352 265674
rect 491300 265610 491352 265616
rect 490012 25560 490064 25566
rect 490012 25502 490064 25508
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 25502
rect 491312 16574 491340 265610
rect 492680 246356 492732 246362
rect 492680 246298 492732 246304
rect 492692 16574 492720 246298
rect 494072 16574 494100 318038
rect 498200 316736 498252 316742
rect 498200 316678 498252 316684
rect 495440 264240 495492 264246
rect 495440 264182 495492 264188
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 264182
rect 496820 243568 496872 243574
rect 496820 243510 496872 243516
rect 496832 16574 496860 243510
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 316678
rect 498292 262880 498344 262886
rect 498292 262822 498344 262828
rect 498304 16574 498332 262822
rect 499580 242208 499632 242214
rect 499580 242150 499632 242156
rect 499592 16574 499620 242150
rect 500972 16574 501000 331910
rect 507860 329112 507912 329118
rect 507860 329054 507912 329060
rect 505100 305652 505152 305658
rect 505100 305594 505152 305600
rect 502340 261520 502392 261526
rect 502340 261462 502392 261468
rect 502352 16574 502380 261462
rect 503720 240780 503772 240786
rect 503720 240722 503772 240728
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 240722
rect 505112 16574 505140 305594
rect 506480 283620 506532 283626
rect 506480 283562 506532 283568
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 283562
rect 506572 26920 506624 26926
rect 506572 26862 506624 26868
rect 506584 16574 506612 26862
rect 507872 16574 507900 329054
rect 514760 327752 514812 327758
rect 514760 327694 514812 327700
rect 512000 313948 512052 313954
rect 512000 313890 512052 313896
rect 509240 260160 509292 260166
rect 509240 260102 509292 260108
rect 509252 16574 509280 260102
rect 510620 239420 510672 239426
rect 510620 239362 510672 239368
rect 510632 16574 510660 239362
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 313890
rect 513380 301504 513432 301510
rect 513380 301446 513432 301452
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 301446
rect 514772 3534 514800 327694
rect 525800 323604 525852 323610
rect 525800 323546 525852 323552
rect 518900 315308 518952 315314
rect 518900 315250 518952 315256
rect 516140 257372 516192 257378
rect 516140 257314 516192 257320
rect 514852 28280 514904 28286
rect 514852 28222 514904 28228
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 28222
rect 516152 16574 516180 257314
rect 517520 238060 517572 238066
rect 517520 238002 517572 238008
rect 517532 16574 517560 238002
rect 518912 16574 518940 315250
rect 520280 282192 520332 282198
rect 520280 282134 520332 282140
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 282134
rect 521660 236700 521712 236706
rect 521660 236642 521712 236648
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 236642
rect 524420 235272 524472 235278
rect 524420 235214 524472 235220
rect 523040 21412 523092 21418
rect 523040 21354 523092 21360
rect 523052 3534 523080 21354
rect 524432 16574 524460 235214
rect 525812 16574 525840 323546
rect 529940 322244 529992 322250
rect 529940 322186 529992 322192
rect 527180 300144 527232 300150
rect 527180 300086 527232 300092
rect 527192 16574 527220 300086
rect 528560 233912 528612 233918
rect 528560 233854 528612 233860
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523132 11756 523184 11762
rect 523132 11698 523184 11704
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 11698
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 233854
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 322186
rect 532700 311160 532752 311166
rect 532700 311102 532752 311108
rect 531320 291848 531372 291854
rect 531320 291790 531372 291796
rect 531332 480 531360 291790
rect 531412 42084 531464 42090
rect 531412 42026 531464 42032
rect 531424 16574 531452 42026
rect 532712 16574 532740 311102
rect 536840 297424 536892 297430
rect 536840 297366 536892 297372
rect 534080 256012 534132 256018
rect 534080 255954 534132 255960
rect 534092 16574 534120 255954
rect 535460 32428 535512 32434
rect 535460 32370 535512 32376
rect 535472 16574 535500 32370
rect 536852 16574 536880 297366
rect 538220 254584 538272 254590
rect 538220 254526 538272 254532
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 254526
rect 539600 231124 539652 231130
rect 539600 231066 539652 231072
rect 539612 480 539640 231066
rect 542360 229764 542412 229770
rect 542360 229706 542412 229712
rect 540980 222896 541032 222902
rect 540980 222838 541032 222844
rect 540992 16574 541020 222838
rect 542372 16574 542400 229706
rect 543752 16574 543780 334562
rect 561680 333260 561732 333266
rect 561680 333202 561732 333208
rect 546500 331900 546552 331906
rect 546500 331842 546552 331848
rect 545120 290488 545172 290494
rect 545120 290430 545172 290436
rect 545132 16574 545160 290430
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540796 4820 540848 4826
rect 540796 4762 540848 4768
rect 540808 480 540836 4762
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 331842
rect 550640 330540 550692 330546
rect 550640 330482 550692 330488
rect 547880 295996 547932 296002
rect 547880 295938 547932 295944
rect 547892 480 547920 295938
rect 547972 253224 548024 253230
rect 547972 253166 548024 253172
rect 547984 16574 548012 253166
rect 550652 16574 550680 330482
rect 554780 309800 554832 309806
rect 554780 309742 554832 309748
rect 552020 280832 552072 280838
rect 552020 280774 552072 280780
rect 552032 16574 552060 280774
rect 553400 228404 553452 228410
rect 553400 228346 553452 228352
rect 553412 16574 553440 228346
rect 547984 16546 548656 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550272 15904 550324 15910
rect 550272 15846 550324 15852
rect 550284 480 550312 15846
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 309742
rect 557540 294636 557592 294642
rect 557540 294578 557592 294584
rect 556160 289128 556212 289134
rect 556160 289070 556212 289076
rect 556172 480 556200 289070
rect 556252 17264 556304 17270
rect 556252 17206 556304 17212
rect 556264 16574 556292 17206
rect 557552 16574 557580 294578
rect 560300 227044 560352 227050
rect 560300 226986 560352 226992
rect 560312 16574 560340 226986
rect 561692 16574 561720 333202
rect 576124 320884 576176 320890
rect 576124 320826 576176 320832
rect 564440 308440 564492 308446
rect 564440 308382 564492 308388
rect 563060 251864 563112 251870
rect 563060 251806 563112 251812
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 559288 13116 559340 13122
rect 559288 13058 559340 13064
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 13058
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 251806
rect 564452 3534 564480 308382
rect 568580 307080 568632 307086
rect 568580 307022 568632 307028
rect 565820 250504 565872 250510
rect 565820 250446 565872 250452
rect 564532 29640 564584 29646
rect 564532 29582 564584 29588
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 29582
rect 565832 16574 565860 250446
rect 567200 225616 567252 225622
rect 567200 225558 567252 225564
rect 567212 16574 567240 225558
rect 568592 16574 568620 307022
rect 572812 293276 572864 293282
rect 572812 293218 572864 293224
rect 571984 287700 572036 287706
rect 571984 287642 572036 287648
rect 569960 249076 570012 249082
rect 569960 249018 570012 249024
rect 569972 16574 570000 249018
rect 571340 36576 571392 36582
rect 571340 36518 571392 36524
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 36518
rect 571996 3058 572024 287642
rect 572824 6914 572852 293218
rect 574100 224256 574152 224262
rect 574100 224198 574152 224204
rect 574112 16574 574140 224198
rect 574112 16546 575152 16574
rect 572732 6886 572852 6914
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 6886
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 16546
rect 576136 3806 576164 320826
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 579712 100700 579764 100706
rect 579712 100642 579764 100648
rect 579724 99521 579752 100642
rect 579710 99512 579766 99521
rect 579710 99447 579766 99456
rect 579988 86964 580040 86970
rect 579988 86906 580040 86912
rect 580000 86193 580028 86906
rect 579986 86184 580042 86193
rect 579986 86119 580042 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 579804 60716 579856 60722
rect 579804 60658 579856 60664
rect 579816 59673 579844 60658
rect 579802 59664 579858 59673
rect 579802 59599 579858 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576124 3800 576176 3806
rect 576124 3742 576176 3748
rect 576320 480 576348 6122
rect 577424 480 577452 8910
rect 580276 6633 580304 458254
rect 580354 326360 580410 326369
rect 580354 326295 580410 326304
rect 580368 33153 580396 326295
rect 580446 302832 580502 302841
rect 580446 302767 580502 302776
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 580460 19825 580488 302767
rect 580446 19816 580502 19825
rect 580446 19751 580502 19760
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 578608 3800 578660 3806
rect 578608 3742 578660 3748
rect 578620 480 578648 3742
rect 581000 3596 581052 3602
rect 581000 3538 581052 3544
rect 581012 480 581040 3538
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 619112 3386 619168
rect 3330 606056 3386 606112
rect 3054 566888 3110 566944
rect 3330 553832 3386 553888
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632032 3570 632088
rect 3606 579944 3662 580000
rect 3698 527856 3754 527912
rect 3882 475632 3938 475688
rect 3514 462576 3570 462632
rect 3422 460128 3478 460184
rect 3330 449520 3386 449576
rect 2962 410488 3018 410544
rect 3514 423544 3570 423600
rect 3422 397432 3478 397488
rect 3238 371320 3294 371376
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 3514 337320 3570 337376
rect 3422 319232 3478 319288
rect 3422 313928 3478 313984
rect 3330 306176 3386 306232
rect 2870 293120 2926 293176
rect 3238 267144 3294 267200
rect 3330 254088 3386 254144
rect 3238 241032 3294 241088
rect 2778 214956 2780 214976
rect 2780 214956 2832 214976
rect 2832 214956 2834 214976
rect 2778 214920 2834 214956
rect 3330 201864 3386 201920
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3330 149776 3386 149832
rect 3054 58520 3110 58576
rect 3606 316648 3662 316704
rect 3606 136720 3662 136776
rect 3514 110608 3570 110664
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3422 45464 3478 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 40038 460264 40094 460320
rect 7562 334600 7618 334656
rect 8942 333240 8998 333296
rect 10322 320728 10378 320784
rect 11794 318008 11850 318064
rect 10414 293120 10470 293176
rect 6458 3304 6514 3360
rect 13082 315288 13138 315344
rect 14462 311072 14518 311128
rect 17222 298696 17278 298752
rect 18694 297336 18750 297392
rect 15934 3440 15990 3496
rect 21362 295976 21418 296032
rect 22742 294480 22798 294536
rect 272016 458224 272072 458280
rect 344374 460264 344430 460320
rect 349158 460128 349214 460184
rect 407578 459720 407634 459776
rect 237654 457408 237710 457464
rect 239218 457408 239274 457464
rect 242346 457408 242402 457464
rect 243910 457408 243966 457464
rect 246670 457408 246726 457464
rect 248234 457408 248290 457464
rect 250258 457408 250314 457464
rect 251822 457408 251878 457464
rect 253386 457408 253442 457464
rect 256514 457408 256570 457464
rect 257710 457408 257766 457464
rect 259274 457408 259330 457464
rect 261298 457408 261354 457464
rect 262862 457408 262918 457464
rect 264518 457408 264574 457464
rect 266082 457408 266138 457464
rect 267554 457408 267610 457464
rect 268750 457408 268806 457464
rect 270590 457408 270646 457464
rect 383842 457408 383898 457464
rect 385406 457408 385462 457464
rect 388626 457408 388682 457464
rect 390190 457408 390246 457464
rect 393502 457408 393558 457464
rect 394882 457408 394938 457464
rect 398102 457408 398158 457464
rect 399666 457408 399722 457464
rect 401230 457408 401286 457464
rect 402978 457408 403034 457464
rect 404358 457408 404414 457464
rect 406014 457408 406070 457464
rect 409142 457408 409198 457464
rect 410706 457408 410762 457464
rect 412270 457408 412326 457464
rect 232594 319368 232650 319424
rect 236182 3304 236238 3360
rect 238758 3440 238814 3496
rect 277122 3304 277178 3360
rect 320270 3304 320326 3360
rect 383014 336776 383070 336832
rect 382278 3440 382334 3496
rect 414202 3304 414258 3360
rect 420182 331744 420238 331800
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 423034 329024 423090 329080
rect 424322 327664 424378 327720
rect 425702 323584 425758 323640
rect 424322 291760 424378 291816
rect 438122 322088 438178 322144
rect 427082 309712 427138 309768
rect 428462 308352 428518 308408
rect 429842 306992 429898 307048
rect 431222 301416 431278 301472
rect 432602 300056 432658 300112
rect 435362 290400 435418 290456
rect 436742 289040 436798 289096
rect 445022 287680 445078 287736
rect 460202 304136 460258 304192
rect 479522 330384 479578 330440
rect 479338 3440 479394 3496
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579618 125976 579674 126032
rect 580170 112784 580226 112840
rect 579710 99456 579766 99512
rect 579986 86128 580042 86184
rect 580170 72936 580226 72992
rect 579802 59608 579858 59664
rect 580170 46280 580226 46336
rect 580354 326304 580410 326360
rect 580446 302776 580502 302832
rect 580354 33088 580410 33144
rect 580446 19760 580502 19816
rect 580262 6568 580318 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3601 580002 3667 580005
rect -960 580000 3667 580002
rect -960 579944 3606 580000
rect 3662 579944 3667 580000
rect -960 579942 3667 579944
rect -960 579852 480 579942
rect 3601 579939 3667 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3693 527914 3759 527917
rect -960 527912 3759 527914
rect -960 527856 3698 527912
rect 3754 527856 3759 527912
rect -960 527854 3759 527856
rect -960 527764 480 527854
rect 3693 527851 3759 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 40033 460322 40099 460325
rect 344369 460322 344435 460325
rect 40033 460320 344435 460322
rect 40033 460264 40038 460320
rect 40094 460264 344374 460320
rect 344430 460264 344435 460320
rect 40033 460262 344435 460264
rect 40033 460259 40099 460262
rect 344369 460259 344435 460262
rect 3417 460186 3483 460189
rect 349153 460186 349219 460189
rect 3417 460184 349219 460186
rect 3417 460128 3422 460184
rect 3478 460128 349158 460184
rect 349214 460128 349219 460184
rect 3417 460126 349219 460128
rect 3417 460123 3483 460126
rect 349153 460123 349219 460126
rect 402094 459716 402100 459780
rect 402164 459778 402170 459780
rect 407573 459778 407639 459781
rect 402164 459776 407639 459778
rect 402164 459720 407578 459776
rect 407634 459720 407639 459776
rect 402164 459718 407639 459720
rect 402164 459716 402170 459718
rect 407573 459715 407639 459718
rect 272011 458282 272077 458285
rect 273846 458282 273852 458284
rect 272011 458280 273852 458282
rect 272011 458224 272016 458280
rect 272072 458224 273852 458280
rect 272011 458222 273852 458224
rect 272011 458219 272077 458222
rect 273846 458220 273852 458222
rect 273916 458220 273922 458284
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 237649 457466 237715 457469
rect 237966 457466 237972 457468
rect 237649 457464 237972 457466
rect 237649 457408 237654 457464
rect 237710 457408 237972 457464
rect 237649 457406 237972 457408
rect 237649 457403 237715 457406
rect 237966 457404 237972 457406
rect 238036 457404 238042 457468
rect 239213 457466 239279 457469
rect 240726 457466 240732 457468
rect 239213 457464 240732 457466
rect 239213 457408 239218 457464
rect 239274 457408 240732 457464
rect 239213 457406 240732 457408
rect 239213 457403 239279 457406
rect 240726 457404 240732 457406
rect 240796 457404 240802 457468
rect 242341 457466 242407 457469
rect 242750 457466 242756 457468
rect 242341 457464 242756 457466
rect 242341 457408 242346 457464
rect 242402 457408 242756 457464
rect 242341 457406 242756 457408
rect 242341 457403 242407 457406
rect 242750 457404 242756 457406
rect 242820 457404 242826 457468
rect 243905 457466 243971 457469
rect 244038 457466 244044 457468
rect 243905 457464 244044 457466
rect 243905 457408 243910 457464
rect 243966 457408 244044 457464
rect 243905 457406 244044 457408
rect 243905 457403 243971 457406
rect 244038 457404 244044 457406
rect 244108 457404 244114 457468
rect 246665 457466 246731 457469
rect 248229 457468 248295 457469
rect 246798 457466 246804 457468
rect 246665 457464 246804 457466
rect 246665 457408 246670 457464
rect 246726 457408 246804 457464
rect 246665 457406 246804 457408
rect 246665 457403 246731 457406
rect 246798 457404 246804 457406
rect 246868 457404 246874 457468
rect 248229 457464 248276 457468
rect 248340 457466 248346 457468
rect 250253 457466 250319 457469
rect 251030 457466 251036 457468
rect 248229 457408 248234 457464
rect 248229 457404 248276 457408
rect 248340 457406 248386 457466
rect 250253 457464 251036 457466
rect 250253 457408 250258 457464
rect 250314 457408 251036 457464
rect 250253 457406 251036 457408
rect 248340 457404 248346 457406
rect 248229 457403 248295 457404
rect 250253 457403 250319 457406
rect 251030 457404 251036 457406
rect 251100 457404 251106 457468
rect 251817 457466 251883 457469
rect 252318 457466 252324 457468
rect 251817 457464 252324 457466
rect 251817 457408 251822 457464
rect 251878 457408 252324 457464
rect 251817 457406 252324 457408
rect 251817 457403 251883 457406
rect 252318 457404 252324 457406
rect 252388 457404 252394 457468
rect 253381 457466 253447 457469
rect 256509 457468 256575 457469
rect 253606 457466 253612 457468
rect 253381 457464 253612 457466
rect 253381 457408 253386 457464
rect 253442 457408 253612 457464
rect 253381 457406 253612 457408
rect 253381 457403 253447 457406
rect 253606 457404 253612 457406
rect 253676 457404 253682 457468
rect 256509 457464 256556 457468
rect 256620 457466 256626 457468
rect 257705 457466 257771 457469
rect 259269 457468 259335 457469
rect 257838 457466 257844 457468
rect 256509 457408 256514 457464
rect 256509 457404 256556 457408
rect 256620 457406 256666 457466
rect 257705 457464 257844 457466
rect 257705 457408 257710 457464
rect 257766 457408 257844 457464
rect 257705 457406 257844 457408
rect 256620 457404 256626 457406
rect 256509 457403 256575 457404
rect 257705 457403 257771 457406
rect 257838 457404 257844 457406
rect 257908 457404 257914 457468
rect 259269 457464 259316 457468
rect 259380 457466 259386 457468
rect 261293 457466 261359 457469
rect 262070 457466 262076 457468
rect 259269 457408 259274 457464
rect 259269 457404 259316 457408
rect 259380 457406 259426 457466
rect 261293 457464 262076 457466
rect 261293 457408 261298 457464
rect 261354 457408 262076 457464
rect 261293 457406 262076 457408
rect 259380 457404 259386 457406
rect 259269 457403 259335 457404
rect 261293 457403 261359 457406
rect 262070 457404 262076 457406
rect 262140 457404 262146 457468
rect 262857 457466 262923 457469
rect 263358 457466 263364 457468
rect 262857 457464 263364 457466
rect 262857 457408 262862 457464
rect 262918 457408 263364 457464
rect 262857 457406 263364 457408
rect 262857 457403 262923 457406
rect 263358 457404 263364 457406
rect 263428 457404 263434 457468
rect 264513 457466 264579 457469
rect 266077 457468 266143 457469
rect 267549 457468 267615 457469
rect 264830 457466 264836 457468
rect 264513 457464 264836 457466
rect 264513 457408 264518 457464
rect 264574 457408 264836 457464
rect 264513 457406 264836 457408
rect 264513 457403 264579 457406
rect 264830 457404 264836 457406
rect 264900 457404 264906 457468
rect 266077 457464 266124 457468
rect 266188 457466 266194 457468
rect 266077 457408 266082 457464
rect 266077 457404 266124 457408
rect 266188 457406 266234 457466
rect 267549 457464 267596 457468
rect 267660 457466 267666 457468
rect 268745 457466 268811 457469
rect 268878 457466 268884 457468
rect 267549 457408 267554 457464
rect 266188 457404 266194 457406
rect 267549 457404 267596 457408
rect 267660 457406 267706 457466
rect 268745 457464 268884 457466
rect 268745 457408 268750 457464
rect 268806 457408 268884 457464
rect 268745 457406 268884 457408
rect 267660 457404 267666 457406
rect 266077 457403 266143 457404
rect 267549 457403 267615 457404
rect 268745 457403 268811 457406
rect 268878 457404 268884 457406
rect 268948 457404 268954 457468
rect 270585 457466 270651 457469
rect 271086 457466 271092 457468
rect 270585 457464 271092 457466
rect 270585 457408 270590 457464
rect 270646 457408 271092 457464
rect 270585 457406 271092 457408
rect 270585 457403 270651 457406
rect 271086 457404 271092 457406
rect 271156 457404 271162 457468
rect 383694 457404 383700 457468
rect 383764 457466 383770 457468
rect 383837 457466 383903 457469
rect 383764 457464 383903 457466
rect 383764 457408 383842 457464
rect 383898 457408 383903 457464
rect 383764 457406 383903 457408
rect 383764 457404 383770 457406
rect 383837 457403 383903 457406
rect 384982 457404 384988 457468
rect 385052 457466 385058 457468
rect 385401 457466 385467 457469
rect 385052 457464 385467 457466
rect 385052 457408 385406 457464
rect 385462 457408 385467 457464
rect 385052 457406 385467 457408
rect 385052 457404 385058 457406
rect 385401 457403 385467 457406
rect 387742 457404 387748 457468
rect 387812 457466 387818 457468
rect 388621 457466 388687 457469
rect 387812 457464 388687 457466
rect 387812 457408 388626 457464
rect 388682 457408 388687 457464
rect 387812 457406 388687 457408
rect 387812 457404 387818 457406
rect 388621 457403 388687 457406
rect 389214 457404 389220 457468
rect 389284 457466 389290 457468
rect 390185 457466 390251 457469
rect 393497 457468 393563 457469
rect 393446 457466 393452 457468
rect 389284 457464 390251 457466
rect 389284 457408 390190 457464
rect 390246 457408 390251 457464
rect 389284 457406 390251 457408
rect 393406 457406 393452 457466
rect 393516 457464 393563 457468
rect 393558 457408 393563 457464
rect 389284 457404 389290 457406
rect 390185 457403 390251 457406
rect 393446 457404 393452 457406
rect 393516 457404 393563 457408
rect 394734 457404 394740 457468
rect 394804 457466 394810 457468
rect 394877 457466 394943 457469
rect 394804 457464 394943 457466
rect 394804 457408 394882 457464
rect 394938 457408 394943 457464
rect 394804 457406 394943 457408
rect 394804 457404 394810 457406
rect 393497 457403 393563 457404
rect 394877 457403 394943 457406
rect 396574 457404 396580 457468
rect 396644 457466 396650 457468
rect 398097 457466 398163 457469
rect 396644 457464 398163 457466
rect 396644 457408 398102 457464
rect 398158 457408 398163 457464
rect 396644 457406 398163 457408
rect 396644 457404 396650 457406
rect 398097 457403 398163 457406
rect 398782 457404 398788 457468
rect 398852 457466 398858 457468
rect 399661 457466 399727 457469
rect 398852 457464 399727 457466
rect 398852 457408 399666 457464
rect 399722 457408 399727 457464
rect 398852 457406 399727 457408
rect 398852 457404 398858 457406
rect 399661 457403 399727 457406
rect 400254 457404 400260 457468
rect 400324 457466 400330 457468
rect 401225 457466 401291 457469
rect 400324 457464 401291 457466
rect 400324 457408 401230 457464
rect 401286 457408 401291 457464
rect 400324 457406 401291 457408
rect 400324 457404 400330 457406
rect 401225 457403 401291 457406
rect 402973 457468 403039 457469
rect 404353 457468 404419 457469
rect 402973 457464 403020 457468
rect 403084 457466 403090 457468
rect 404302 457466 404308 457468
rect 402973 457408 402978 457464
rect 402973 457404 403020 457408
rect 403084 457406 403130 457466
rect 404262 457406 404308 457466
rect 404372 457464 404419 457468
rect 404414 457408 404419 457464
rect 403084 457404 403090 457406
rect 404302 457404 404308 457406
rect 404372 457404 404419 457408
rect 405774 457404 405780 457468
rect 405844 457466 405850 457468
rect 406009 457466 406075 457469
rect 405844 457464 406075 457466
rect 405844 457408 406014 457464
rect 406070 457408 406075 457464
rect 405844 457406 406075 457408
rect 405844 457404 405850 457406
rect 402973 457403 403039 457404
rect 404353 457403 404419 457404
rect 406009 457403 406075 457406
rect 408718 457404 408724 457468
rect 408788 457466 408794 457468
rect 409137 457466 409203 457469
rect 408788 457464 409203 457466
rect 408788 457408 409142 457464
rect 409198 457408 409203 457464
rect 408788 457406 409203 457408
rect 408788 457404 408794 457406
rect 409137 457403 409203 457406
rect 409822 457404 409828 457468
rect 409892 457466 409898 457468
rect 410701 457466 410767 457469
rect 409892 457464 410767 457466
rect 409892 457408 410706 457464
rect 410762 457408 410767 457464
rect 409892 457406 410767 457408
rect 409892 457404 409898 457406
rect 410701 457403 410767 457406
rect 411294 457404 411300 457468
rect 411364 457466 411370 457468
rect 412265 457466 412331 457469
rect 411364 457464 412331 457466
rect 411364 457408 412270 457464
rect 412326 457408 412331 457464
rect 411364 457406 412331 457408
rect 411364 457404 411370 457406
rect 412265 457403 412331 457406
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect 3509 337378 3575 337381
rect 400254 337378 400260 337380
rect 3509 337376 400260 337378
rect 3509 337320 3514 337376
rect 3570 337320 400260 337376
rect 3509 337318 400260 337320
rect 3509 337315 3575 337318
rect 400254 337316 400260 337318
rect 400324 337316 400330 337380
rect 383009 336834 383075 336837
rect 384982 336834 384988 336836
rect 383009 336832 384988 336834
rect 383009 336776 383014 336832
rect 383070 336776 384988 336832
rect 383009 336774 384988 336776
rect 383009 336771 383075 336774
rect 384982 336772 384988 336774
rect 385052 336772 385058 336836
rect 7557 334658 7623 334661
rect 405774 334658 405780 334660
rect 7557 334656 405780 334658
rect 7557 334600 7562 334656
rect 7618 334600 405780 334656
rect 7557 334598 405780 334600
rect 7557 334595 7623 334598
rect 405774 334596 405780 334598
rect 405844 334596 405850 334660
rect 8937 333298 9003 333301
rect 409822 333298 409828 333300
rect 8937 333296 409828 333298
rect 8937 333240 8942 333296
rect 8998 333240 409828 333296
rect 8937 333238 409828 333240
rect 8937 333235 9003 333238
rect 409822 333236 409828 333238
rect 409892 333236 409898 333300
rect -960 332196 480 332436
rect 251030 331740 251036 331804
rect 251100 331802 251106 331804
rect 420177 331802 420243 331805
rect 251100 331800 420243 331802
rect 251100 331744 420182 331800
rect 420238 331744 420243 331800
rect 251100 331742 420243 331744
rect 251100 331740 251106 331742
rect 420177 331739 420243 331742
rect 259310 330380 259316 330444
rect 259380 330442 259386 330444
rect 479517 330442 479583 330445
rect 259380 330440 479583 330442
rect 259380 330384 479522 330440
rect 479578 330384 479583 330440
rect 259380 330382 479583 330384
rect 259380 330380 259386 330382
rect 479517 330379 479583 330382
rect 264830 329020 264836 329084
rect 264900 329082 264906 329084
rect 423029 329082 423095 329085
rect 264900 329080 423095 329082
rect 264900 329024 423034 329080
rect 423090 329024 423095 329080
rect 264900 329022 423095 329024
rect 264900 329020 264906 329022
rect 423029 329019 423095 329022
rect 268878 327660 268884 327724
rect 268948 327722 268954 327724
rect 424317 327722 424383 327725
rect 268948 327720 424383 327722
rect 268948 327664 424322 327720
rect 424378 327664 424383 327720
rect 268948 327662 424383 327664
rect 268948 327660 268954 327662
rect 424317 327659 424383 327662
rect 237966 326300 237972 326364
rect 238036 326362 238042 326364
rect 580349 326362 580415 326365
rect 238036 326360 580415 326362
rect 238036 326304 580354 326360
rect 580410 326304 580415 326360
rect 238036 326302 580415 326304
rect 238036 326300 238042 326302
rect 580349 326299 580415 326302
rect 583520 325274 584960 325364
rect 583342 325214 584960 325274
rect 583342 325138 583402 325214
rect 583520 325138 584960 325214
rect 583342 325124 584960 325138
rect 583342 325078 583586 325124
rect 271086 324396 271092 324460
rect 271156 324458 271162 324460
rect 583526 324458 583586 325078
rect 271156 324398 583586 324458
rect 271156 324396 271162 324398
rect 242750 323580 242756 323644
rect 242820 323642 242826 323644
rect 425697 323642 425763 323645
rect 242820 323640 425763 323642
rect 242820 323584 425702 323640
rect 425758 323584 425763 323640
rect 242820 323582 425763 323584
rect 242820 323580 242826 323582
rect 425697 323579 425763 323582
rect 246798 322084 246804 322148
rect 246868 322146 246874 322148
rect 438117 322146 438183 322149
rect 246868 322144 438183 322146
rect 246868 322088 438122 322144
rect 438178 322088 438183 322144
rect 246868 322086 438183 322088
rect 246868 322084 246874 322086
rect 438117 322083 438183 322086
rect 10317 320786 10383 320789
rect 383694 320786 383700 320788
rect 10317 320784 383700 320786
rect 10317 320728 10322 320784
rect 10378 320728 383700 320784
rect 10317 320726 383700 320728
rect 10317 320723 10383 320726
rect 383694 320724 383700 320726
rect 383764 320724 383770 320788
rect 232589 319426 232655 319429
rect 387742 319426 387748 319428
rect 232589 319424 387748 319426
rect -960 319290 480 319380
rect 232589 319368 232594 319424
rect 232650 319368 387748 319424
rect 232589 319366 387748 319368
rect 232589 319363 232655 319366
rect 387742 319364 387748 319366
rect 387812 319364 387818 319428
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 11789 318066 11855 318069
rect 393078 318066 393084 318068
rect 11789 318064 393084 318066
rect 11789 318008 11794 318064
rect 11850 318008 393084 318064
rect 11789 318006 393084 318008
rect 11789 318003 11855 318006
rect 393078 318004 393084 318006
rect 393148 318004 393154 318068
rect 3601 316706 3667 316709
rect 396574 316706 396580 316708
rect 3601 316704 396580 316706
rect 3601 316648 3606 316704
rect 3662 316648 396580 316704
rect 3601 316646 396580 316648
rect 3601 316643 3667 316646
rect 396574 316644 396580 316646
rect 396644 316644 396650 316708
rect 13077 315346 13143 315349
rect 403014 315346 403020 315348
rect 13077 315344 403020 315346
rect 13077 315288 13082 315344
rect 13138 315288 403020 315344
rect 13077 315286 403020 315288
rect 13077 315283 13143 315286
rect 403014 315284 403020 315286
rect 403084 315284 403090 315348
rect 3417 313986 3483 313989
rect 402094 313986 402100 313988
rect 3417 313984 402100 313986
rect 3417 313928 3422 313984
rect 3478 313928 402100 313984
rect 3417 313926 402100 313928
rect 3417 313923 3483 313926
rect 402094 313924 402100 313926
rect 402164 313924 402170 313988
rect 583520 312082 584960 312172
rect 567150 312022 584960 312082
rect 273846 311884 273852 311948
rect 273916 311946 273922 311948
rect 567150 311946 567210 312022
rect 273916 311886 567210 311946
rect 583520 311932 584960 312022
rect 273916 311884 273922 311886
rect 14457 311130 14523 311133
rect 411294 311130 411300 311132
rect 14457 311128 411300 311130
rect 14457 311072 14462 311128
rect 14518 311072 411300 311128
rect 14457 311070 411300 311072
rect 14457 311067 14523 311070
rect 411294 311068 411300 311070
rect 411364 311068 411370 311132
rect 252318 309708 252324 309772
rect 252388 309770 252394 309772
rect 427077 309770 427143 309773
rect 252388 309768 427143 309770
rect 252388 309712 427082 309768
rect 427138 309712 427143 309768
rect 252388 309710 427143 309712
rect 252388 309708 252394 309710
rect 427077 309707 427143 309710
rect 256550 308348 256556 308412
rect 256620 308410 256626 308412
rect 428457 308410 428523 308413
rect 256620 308408 428523 308410
rect 256620 308352 428462 308408
rect 428518 308352 428523 308408
rect 256620 308350 428523 308352
rect 256620 308348 256626 308350
rect 428457 308347 428523 308350
rect 262070 306988 262076 307052
rect 262140 307050 262146 307052
rect 429837 307050 429903 307053
rect 262140 307048 429903 307050
rect 262140 306992 429842 307048
rect 429898 306992 429903 307048
rect 262140 306990 429903 306992
rect 262140 306988 262146 306990
rect 429837 306987 429903 306990
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 266118 304132 266124 304196
rect 266188 304194 266194 304196
rect 460197 304194 460263 304197
rect 266188 304192 460263 304194
rect 266188 304136 460202 304192
rect 460258 304136 460263 304192
rect 266188 304134 460263 304136
rect 266188 304132 266194 304134
rect 460197 304131 460263 304134
rect 240726 302772 240732 302836
rect 240796 302834 240802 302836
rect 580441 302834 580507 302837
rect 240796 302832 580507 302834
rect 240796 302776 580446 302832
rect 580502 302776 580507 302832
rect 240796 302774 580507 302776
rect 240796 302772 240802 302774
rect 580441 302771 580507 302774
rect 244038 301412 244044 301476
rect 244108 301474 244114 301476
rect 431217 301474 431283 301477
rect 244108 301472 431283 301474
rect 244108 301416 431222 301472
rect 431278 301416 431283 301472
rect 244108 301414 431283 301416
rect 244108 301412 244114 301414
rect 431217 301411 431283 301414
rect 248270 300052 248276 300116
rect 248340 300114 248346 300116
rect 432597 300114 432663 300117
rect 248340 300112 432663 300114
rect 248340 300056 432602 300112
rect 432658 300056 432663 300112
rect 248340 300054 432663 300056
rect 248340 300052 248346 300054
rect 432597 300051 432663 300054
rect 17217 298754 17283 298757
rect 389214 298754 389220 298756
rect 17217 298752 389220 298754
rect 17217 298696 17222 298752
rect 17278 298696 389220 298752
rect 17217 298694 389220 298696
rect 17217 298691 17283 298694
rect 389214 298692 389220 298694
rect 389284 298692 389290 298756
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 18689 297394 18755 297397
rect 394734 297394 394740 297396
rect 18689 297392 394740 297394
rect 18689 297336 18694 297392
rect 18750 297336 394740 297392
rect 18689 297334 394740 297336
rect 18689 297331 18755 297334
rect 394734 297332 394740 297334
rect 394804 297332 394810 297396
rect 21357 296034 21423 296037
rect 398782 296034 398788 296036
rect 21357 296032 398788 296034
rect 21357 295976 21362 296032
rect 21418 295976 398788 296032
rect 21357 295974 398788 295976
rect 21357 295971 21423 295974
rect 398782 295972 398788 295974
rect 398852 295972 398858 296036
rect 22737 294538 22803 294541
rect 404302 294538 404308 294540
rect 22737 294536 404308 294538
rect 22737 294480 22742 294536
rect 22798 294480 404308 294536
rect 22737 294478 404308 294480
rect 22737 294475 22803 294478
rect 404302 294476 404308 294478
rect 404372 294476 404378 294540
rect -960 293178 480 293268
rect 2865 293178 2931 293181
rect -960 293176 2931 293178
rect -960 293120 2870 293176
rect 2926 293120 2931 293176
rect -960 293118 2931 293120
rect -960 293028 480 293118
rect 2865 293115 2931 293118
rect 10409 293178 10475 293181
rect 408718 293178 408724 293180
rect 10409 293176 408724 293178
rect 10409 293120 10414 293176
rect 10470 293120 408724 293176
rect 10409 293118 408724 293120
rect 10409 293115 10475 293118
rect 408718 293116 408724 293118
rect 408788 293116 408794 293180
rect 253606 291756 253612 291820
rect 253676 291818 253682 291820
rect 424317 291818 424383 291821
rect 253676 291816 424383 291818
rect 253676 291760 424322 291816
rect 424378 291760 424383 291816
rect 253676 291758 424383 291760
rect 253676 291756 253682 291758
rect 424317 291755 424383 291758
rect 257838 290396 257844 290460
rect 257908 290458 257914 290460
rect 435357 290458 435423 290461
rect 257908 290456 435423 290458
rect 257908 290400 435362 290456
rect 435418 290400 435423 290456
rect 257908 290398 435423 290400
rect 257908 290396 257914 290398
rect 435357 290395 435423 290398
rect 263358 289036 263364 289100
rect 263428 289098 263434 289100
rect 436737 289098 436803 289101
rect 263428 289096 436803 289098
rect 263428 289040 436742 289096
rect 436798 289040 436803 289096
rect 263428 289038 436803 289040
rect 263428 289036 263434 289038
rect 436737 289035 436803 289038
rect 267590 287676 267596 287740
rect 267660 287738 267666 287740
rect 445017 287738 445083 287741
rect 267660 287736 445083 287738
rect 267660 287680 445022 287736
rect 445078 287680 445083 287736
rect 267660 287678 445083 287680
rect 267660 287676 267666 287678
rect 445017 287675 445083 287678
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3509 110666 3575 110669
rect -960 110664 3575 110666
rect -960 110608 3514 110664
rect 3570 110608 3575 110664
rect -960 110606 3575 110608
rect -960 110516 480 110606
rect 3509 110603 3575 110606
rect 579705 99514 579771 99517
rect 583520 99514 584960 99604
rect 579705 99512 584960 99514
rect 579705 99456 579710 99512
rect 579766 99456 584960 99512
rect 579705 99454 584960 99456
rect 579705 99451 579771 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 579981 86186 580047 86189
rect 583520 86186 584960 86276
rect 579981 86184 584960 86186
rect 579981 86128 579986 86184
rect 580042 86128 584960 86184
rect 579981 86126 584960 86128
rect 579981 86123 580047 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 579797 59666 579863 59669
rect 583520 59666 584960 59756
rect 579797 59664 584960 59666
rect 579797 59608 579802 59664
rect 579858 59608 584960 59664
rect 579797 59606 584960 59608
rect 579797 59603 579863 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 580441 19818 580507 19821
rect 583520 19818 584960 19908
rect 580441 19816 584960 19818
rect 580441 19760 580446 19816
rect 580502 19760 584960 19816
rect 580441 19758 584960 19760
rect 580441 19755 580507 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 15929 3498 15995 3501
rect 238753 3498 238819 3501
rect 15929 3496 238819 3498
rect 15929 3440 15934 3496
rect 15990 3440 238758 3496
rect 238814 3440 238819 3496
rect 15929 3438 238819 3440
rect 15929 3435 15995 3438
rect 238753 3435 238819 3438
rect 382273 3498 382339 3501
rect 479333 3498 479399 3501
rect 382273 3496 479399 3498
rect 382273 3440 382278 3496
rect 382334 3440 479338 3496
rect 479394 3440 479399 3496
rect 382273 3438 479399 3440
rect 382273 3435 382339 3438
rect 479333 3435 479399 3438
rect 6453 3362 6519 3365
rect 236177 3362 236243 3365
rect 6453 3360 236243 3362
rect 6453 3304 6458 3360
rect 6514 3304 236182 3360
rect 236238 3304 236243 3360
rect 6453 3302 236243 3304
rect 6453 3299 6519 3302
rect 236177 3299 236243 3302
rect 277117 3362 277183 3365
rect 320265 3362 320331 3365
rect 277117 3360 320331 3362
rect 277117 3304 277122 3360
rect 277178 3304 320270 3360
rect 320326 3304 320331 3360
rect 277117 3302 320331 3304
rect 277117 3299 277183 3302
rect 320265 3299 320331 3302
rect 414197 3362 414263 3365
rect 583385 3362 583451 3365
rect 414197 3360 583451 3362
rect 414197 3304 414202 3360
rect 414258 3304 583390 3360
rect 583446 3304 583451 3360
rect 414197 3302 583451 3304
rect 414197 3299 414263 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 402100 459716 402164 459780
rect 273852 458220 273916 458284
rect 237972 457404 238036 457468
rect 240732 457404 240796 457468
rect 242756 457404 242820 457468
rect 244044 457404 244108 457468
rect 246804 457404 246868 457468
rect 248276 457464 248340 457468
rect 248276 457408 248290 457464
rect 248290 457408 248340 457464
rect 248276 457404 248340 457408
rect 251036 457404 251100 457468
rect 252324 457404 252388 457468
rect 253612 457404 253676 457468
rect 256556 457464 256620 457468
rect 256556 457408 256570 457464
rect 256570 457408 256620 457464
rect 256556 457404 256620 457408
rect 257844 457404 257908 457468
rect 259316 457464 259380 457468
rect 259316 457408 259330 457464
rect 259330 457408 259380 457464
rect 259316 457404 259380 457408
rect 262076 457404 262140 457468
rect 263364 457404 263428 457468
rect 264836 457404 264900 457468
rect 266124 457464 266188 457468
rect 266124 457408 266138 457464
rect 266138 457408 266188 457464
rect 266124 457404 266188 457408
rect 267596 457464 267660 457468
rect 267596 457408 267610 457464
rect 267610 457408 267660 457464
rect 267596 457404 267660 457408
rect 268884 457404 268948 457468
rect 271092 457404 271156 457468
rect 383700 457404 383764 457468
rect 384988 457404 385052 457468
rect 387748 457404 387812 457468
rect 389220 457404 389284 457468
rect 393452 457464 393516 457468
rect 393452 457408 393502 457464
rect 393502 457408 393516 457464
rect 393452 457404 393516 457408
rect 394740 457404 394804 457468
rect 396580 457404 396644 457468
rect 398788 457404 398852 457468
rect 400260 457404 400324 457468
rect 403020 457464 403084 457468
rect 403020 457408 403034 457464
rect 403034 457408 403084 457464
rect 403020 457404 403084 457408
rect 404308 457464 404372 457468
rect 404308 457408 404358 457464
rect 404358 457408 404372 457464
rect 404308 457404 404372 457408
rect 405780 457404 405844 457468
rect 408724 457404 408788 457468
rect 409828 457404 409892 457468
rect 411300 457404 411364 457468
rect 400260 337316 400324 337380
rect 384988 336772 385052 336836
rect 405780 334596 405844 334660
rect 409828 333236 409892 333300
rect 251036 331740 251100 331804
rect 259316 330380 259380 330444
rect 264836 329020 264900 329084
rect 268884 327660 268948 327724
rect 237972 326300 238036 326364
rect 271092 324396 271156 324460
rect 242756 323580 242820 323644
rect 246804 322084 246868 322148
rect 383700 320724 383764 320788
rect 387748 319364 387812 319428
rect 393084 318004 393148 318068
rect 396580 316644 396644 316708
rect 403020 315284 403084 315348
rect 402100 313924 402164 313988
rect 273852 311884 273916 311948
rect 411300 311068 411364 311132
rect 252324 309708 252388 309772
rect 256556 308348 256620 308412
rect 262076 306988 262140 307052
rect 266124 304132 266188 304196
rect 240732 302772 240796 302836
rect 244044 301412 244108 301476
rect 248276 300052 248340 300116
rect 389220 298692 389284 298756
rect 394740 297332 394804 297396
rect 398788 295972 398852 296036
rect 404308 294476 404372 294540
rect 408724 293116 408788 293180
rect 253612 291756 253676 291820
rect 257844 290396 257908 290460
rect 263364 289036 263428 289100
rect 267596 287676 267660 287740
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 237971 457468 238037 457469
rect 237971 457404 237972 457468
rect 238036 457404 238037 457468
rect 237971 457403 238037 457404
rect 240731 457468 240797 457469
rect 240731 457404 240732 457468
rect 240796 457404 240797 457468
rect 240731 457403 240797 457404
rect 242755 457468 242821 457469
rect 242755 457404 242756 457468
rect 242820 457404 242821 457468
rect 242755 457403 242821 457404
rect 244043 457468 244109 457469
rect 244043 457404 244044 457468
rect 244108 457404 244109 457468
rect 244043 457403 244109 457404
rect 246803 457468 246869 457469
rect 246803 457404 246804 457468
rect 246868 457404 246869 457468
rect 246803 457403 246869 457404
rect 248275 457468 248341 457469
rect 248275 457404 248276 457468
rect 248340 457404 248341 457468
rect 248275 457403 248341 457404
rect 251035 457468 251101 457469
rect 251035 457404 251036 457468
rect 251100 457404 251101 457468
rect 251035 457403 251101 457404
rect 252323 457468 252389 457469
rect 252323 457404 252324 457468
rect 252388 457404 252389 457468
rect 252323 457403 252389 457404
rect 253611 457468 253677 457469
rect 253611 457404 253612 457468
rect 253676 457404 253677 457468
rect 253611 457403 253677 457404
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 237974 326365 238034 457403
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 237971 326364 238037 326365
rect 237971 326300 237972 326364
rect 238036 326300 238037 326364
rect 237971 326299 238037 326300
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 240734 302837 240794 457403
rect 242758 323645 242818 457403
rect 242755 323644 242821 323645
rect 242755 323580 242756 323644
rect 242820 323580 242821 323644
rect 242755 323579 242821 323580
rect 240731 302836 240797 302837
rect 240731 302772 240732 302836
rect 240796 302772 240797 302836
rect 240731 302771 240797 302772
rect 244046 301477 244106 457403
rect 246806 322149 246866 457403
rect 246803 322148 246869 322149
rect 246803 322084 246804 322148
rect 246868 322084 246869 322148
rect 246803 322083 246869 322084
rect 244043 301476 244109 301477
rect 244043 301412 244044 301476
rect 244108 301412 244109 301476
rect 244043 301411 244109 301412
rect 248278 300117 248338 457403
rect 251038 331805 251098 457403
rect 251035 331804 251101 331805
rect 251035 331740 251036 331804
rect 251100 331740 251101 331804
rect 251035 331739 251101 331740
rect 252326 309773 252386 457403
rect 252323 309772 252389 309773
rect 252323 309708 252324 309772
rect 252388 309708 252389 309772
rect 252323 309707 252389 309708
rect 248275 300116 248341 300117
rect 248275 300052 248276 300116
rect 248340 300052 248341 300116
rect 248275 300051 248341 300052
rect 253614 291821 253674 457403
rect 253794 435454 254414 470898
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 256555 457468 256621 457469
rect 256555 457404 256556 457468
rect 256620 457404 256621 457468
rect 256555 457403 256621 457404
rect 257843 457468 257909 457469
rect 257843 457404 257844 457468
rect 257908 457404 257909 457468
rect 257843 457403 257909 457404
rect 259315 457468 259381 457469
rect 259315 457404 259316 457468
rect 259380 457404 259381 457468
rect 259315 457403 259381 457404
rect 262075 457468 262141 457469
rect 262075 457404 262076 457468
rect 262140 457404 262141 457468
rect 262075 457403 262141 457404
rect 263363 457468 263429 457469
rect 263363 457404 263364 457468
rect 263428 457404 263429 457468
rect 263363 457403 263429 457404
rect 264835 457468 264901 457469
rect 264835 457404 264836 457468
rect 264900 457404 264901 457468
rect 264835 457403 264901 457404
rect 266123 457468 266189 457469
rect 266123 457404 266124 457468
rect 266188 457404 266189 457468
rect 266123 457403 266189 457404
rect 267595 457468 267661 457469
rect 267595 457404 267596 457468
rect 267660 457404 267661 457468
rect 267595 457403 267661 457404
rect 268883 457468 268949 457469
rect 268883 457404 268884 457468
rect 268948 457404 268949 457468
rect 268883 457403 268949 457404
rect 271091 457468 271157 457469
rect 271091 457404 271092 457468
rect 271156 457404 271157 457468
rect 271091 457403 271157 457404
rect 254568 453454 254888 453486
rect 254568 453218 254610 453454
rect 254846 453218 254888 453454
rect 254568 453134 254888 453218
rect 254568 452898 254610 453134
rect 254846 452898 254888 453134
rect 254568 452866 254888 452898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 254568 417454 254888 417486
rect 254568 417218 254610 417454
rect 254846 417218 254888 417454
rect 254568 417134 254888 417218
rect 254568 416898 254610 417134
rect 254846 416898 254888 417134
rect 254568 416866 254888 416898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253611 291820 253677 291821
rect 253611 291756 253612 291820
rect 253676 291756 253677 291820
rect 253611 291755 253677 291756
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 253794 291454 254414 326898
rect 256558 308413 256618 457403
rect 256555 308412 256621 308413
rect 256555 308348 256556 308412
rect 256620 308348 256621 308412
rect 256555 308347 256621 308348
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 257846 290461 257906 457403
rect 259318 330445 259378 457403
rect 259315 330444 259381 330445
rect 259315 330380 259316 330444
rect 259380 330380 259381 330444
rect 259315 330379 259381 330380
rect 262078 307053 262138 457403
rect 262075 307052 262141 307053
rect 262075 306988 262076 307052
rect 262140 306988 262141 307052
rect 262075 306987 262141 306988
rect 257843 290460 257909 290461
rect 257843 290396 257844 290460
rect 257908 290396 257909 290460
rect 257843 290395 257909 290396
rect 263366 289101 263426 457403
rect 264838 329085 264898 457403
rect 264835 329084 264901 329085
rect 264835 329020 264836 329084
rect 264900 329020 264901 329084
rect 264835 329019 264901 329020
rect 266126 304197 266186 457403
rect 266123 304196 266189 304197
rect 266123 304132 266124 304196
rect 266188 304132 266189 304196
rect 266123 304131 266189 304132
rect 263363 289100 263429 289101
rect 263363 289036 263364 289100
rect 263428 289036 263429 289100
rect 263363 289035 263429 289036
rect 267598 287741 267658 457403
rect 268886 327725 268946 457403
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 268883 327724 268949 327725
rect 268883 327660 268884 327724
rect 268948 327660 268949 327724
rect 268883 327659 268949 327660
rect 271094 324461 271154 457403
rect 271794 453454 272414 488898
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 273851 458284 273917 458285
rect 273851 458220 273852 458284
rect 273916 458220 273917 458284
rect 273851 458219 273917 458220
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271091 324460 271157 324461
rect 271091 324396 271092 324460
rect 271156 324396 271157 324460
rect 271091 324395 271157 324396
rect 271794 309454 272414 344898
rect 273854 311949 273914 458219
rect 285288 453454 285608 453486
rect 285288 453218 285330 453454
rect 285566 453218 285608 453454
rect 285288 453134 285608 453218
rect 285288 452898 285330 453134
rect 285566 452898 285608 453134
rect 285288 452866 285608 452898
rect 289794 435454 290414 470898
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 285288 417454 285608 417486
rect 285288 417218 285330 417454
rect 285566 417218 285608 417454
rect 285288 417134 285608 417218
rect 285288 416898 285330 417134
rect 285566 416898 285608 417134
rect 285288 416866 285608 416898
rect 289794 399454 290414 434898
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 307794 417454 308414 452898
rect 316008 453454 316328 453486
rect 316008 453218 316050 453454
rect 316286 453218 316328 453454
rect 316008 453134 316328 453218
rect 316008 452898 316050 453134
rect 316286 452898 316328 453134
rect 316008 452866 316328 452898
rect 325794 435454 326414 470898
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 285288 381454 285608 381486
rect 285288 381218 285330 381454
rect 285566 381218 285608 381454
rect 285288 381134 285608 381218
rect 285288 380898 285330 381134
rect 285566 380898 285608 381134
rect 285288 380866 285608 380898
rect 289794 363454 290414 398898
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 307794 381454 308414 416898
rect 316008 417454 316328 417486
rect 316008 417218 316050 417454
rect 316286 417218 316328 417454
rect 316008 417134 316328 417218
rect 316008 416898 316050 417134
rect 316286 416898 316328 417134
rect 316008 416866 316328 416898
rect 325794 399454 326414 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 343794 417454 344414 452898
rect 346728 453454 347048 453486
rect 346728 453218 346770 453454
rect 347006 453218 347048 453454
rect 346728 453134 347048 453218
rect 346728 452898 346770 453134
rect 347006 452898 347048 453134
rect 346728 452866 347048 452898
rect 361794 435454 362414 470898
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 377448 453454 377768 453486
rect 377448 453218 377490 453454
rect 377726 453218 377768 453454
rect 377448 453134 377768 453218
rect 377448 452898 377490 453134
rect 377726 452898 377768 453134
rect 377448 452866 377768 452898
rect 379794 453454 380414 488898
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 383699 457468 383765 457469
rect 383699 457404 383700 457468
rect 383764 457404 383765 457468
rect 383699 457403 383765 457404
rect 384987 457468 385053 457469
rect 384987 457404 384988 457468
rect 385052 457404 385053 457468
rect 384987 457403 385053 457404
rect 387747 457468 387813 457469
rect 387747 457404 387748 457468
rect 387812 457404 387813 457468
rect 387747 457403 387813 457404
rect 389219 457468 389285 457469
rect 389219 457404 389220 457468
rect 389284 457404 389285 457468
rect 389219 457403 389285 457404
rect 393451 457468 393517 457469
rect 393451 457404 393452 457468
rect 393516 457404 393517 457468
rect 393451 457403 393517 457404
rect 394739 457468 394805 457469
rect 394739 457404 394740 457468
rect 394804 457404 394805 457468
rect 394739 457403 394805 457404
rect 396579 457468 396645 457469
rect 396579 457404 396580 457468
rect 396644 457404 396645 457468
rect 396579 457403 396645 457404
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 361794 435218 361826 435454
rect 362062 435218 362130 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362130 435134
rect 362382 434898 362414 435134
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 289794 327454 290414 362898
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 273851 311948 273917 311949
rect 273851 311884 273852 311948
rect 273916 311884 273917 311948
rect 273851 311883 273917 311884
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 267595 287740 267661 287741
rect 267595 287676 267596 287740
rect 267660 287676 267661 287740
rect 267595 287675 267661 287676
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 307794 345454 308414 380898
rect 316008 381454 316328 381486
rect 316008 381218 316050 381454
rect 316286 381218 316328 381454
rect 316008 381134 316328 381218
rect 316008 380898 316050 381134
rect 316286 380898 316328 381134
rect 316008 380866 316328 380898
rect 325794 363454 326414 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 343794 381454 344414 416898
rect 346728 417454 347048 417486
rect 346728 417218 346770 417454
rect 347006 417218 347048 417454
rect 346728 417134 347048 417218
rect 346728 416898 346770 417134
rect 347006 416898 347048 417134
rect 346728 416866 347048 416898
rect 361794 399454 362414 434898
rect 377448 417454 377768 417486
rect 377448 417218 377490 417454
rect 377726 417218 377768 417454
rect 377448 417134 377768 417218
rect 377448 416898 377490 417134
rect 377726 416898 377768 417134
rect 377448 416866 377768 416898
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 361794 399218 361826 399454
rect 362062 399218 362130 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362130 399134
rect 362382 398898 362414 399134
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 316008 345454 316328 345486
rect 316008 345218 316050 345454
rect 316286 345218 316328 345454
rect 316008 345134 316328 345218
rect 316008 344898 316050 345134
rect 316286 344898 316328 345134
rect 316008 344866 316328 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 325794 327454 326414 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 343794 345454 344414 380898
rect 346728 381454 347048 381486
rect 346728 381218 346770 381454
rect 347006 381218 347048 381454
rect 346728 381134 347048 381218
rect 346728 380898 346770 381134
rect 347006 380898 347048 381134
rect 346728 380866 347048 380898
rect 361794 363454 362414 398898
rect 377448 381454 377768 381486
rect 377448 381218 377490 381454
rect 377726 381218 377768 381454
rect 377448 381134 377768 381218
rect 377448 380898 377490 381134
rect 377726 380898 377768 381134
rect 377448 380866 377768 380898
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 361794 363218 361826 363454
rect 362062 363218 362130 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362130 363134
rect 362382 362898 362414 363134
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 346728 345454 347048 345486
rect 346728 345218 346770 345454
rect 347006 345218 347048 345454
rect 346728 345134 347048 345218
rect 346728 344898 346770 345134
rect 347006 344898 347048 345134
rect 346728 344866 347048 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 361794 327454 362414 362898
rect 377448 345454 377768 345486
rect 377448 345218 377490 345454
rect 377726 345218 377768 345454
rect 377448 345134 377768 345218
rect 377448 344898 377490 345134
rect 377726 344898 377768 345134
rect 377448 344866 377768 344898
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 379794 309454 380414 344898
rect 383702 320789 383762 457403
rect 384990 336837 385050 457403
rect 384987 336836 385053 336837
rect 384987 336772 384988 336836
rect 385052 336772 385053 336836
rect 384987 336771 385053 336772
rect 383699 320788 383765 320789
rect 383699 320724 383700 320788
rect 383764 320724 383765 320788
rect 383699 320723 383765 320724
rect 387750 319429 387810 457403
rect 387747 319428 387813 319429
rect 387747 319364 387748 319428
rect 387812 319364 387813 319428
rect 387747 319363 387813 319364
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 389222 298757 389282 457403
rect 392808 435454 393128 435486
rect 392808 435218 392850 435454
rect 393086 435218 393128 435454
rect 392808 435134 393128 435218
rect 392808 434898 392850 435134
rect 393086 434898 393128 435134
rect 392808 434866 393128 434898
rect 392808 399454 393128 399486
rect 392808 399218 392850 399454
rect 393086 399218 393128 399454
rect 392808 399134 393128 399218
rect 392808 398898 392850 399134
rect 393086 398898 393128 399134
rect 392808 398866 393128 398898
rect 392808 363454 393128 363486
rect 392808 363218 392850 363454
rect 393086 363218 393128 363454
rect 392808 363134 393128 363218
rect 392808 362898 392850 363134
rect 393086 362898 393128 363134
rect 392808 362866 393128 362898
rect 393454 339690 393514 457403
rect 393086 339630 393514 339690
rect 393086 318069 393146 339630
rect 393083 318068 393149 318069
rect 393083 318004 393084 318068
rect 393148 318004 393149 318068
rect 393083 318003 393149 318004
rect 389219 298756 389285 298757
rect 389219 298692 389220 298756
rect 389284 298692 389285 298756
rect 389219 298691 389285 298692
rect 394742 297397 394802 457403
rect 396582 316709 396642 457403
rect 397794 435454 398414 470898
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 402099 459780 402165 459781
rect 402099 459716 402100 459780
rect 402164 459716 402165 459780
rect 402099 459715 402165 459716
rect 398787 457468 398853 457469
rect 398787 457404 398788 457468
rect 398852 457404 398853 457468
rect 398787 457403 398853 457404
rect 400259 457468 400325 457469
rect 400259 457404 400260 457468
rect 400324 457404 400325 457468
rect 400259 457403 400325 457404
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 398790 331230 398850 457403
rect 400262 337381 400322 457403
rect 400259 337380 400325 337381
rect 400259 337316 400260 337380
rect 400324 337316 400325 337380
rect 400259 337315 400325 337316
rect 398790 331170 399034 331230
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 396579 316708 396645 316709
rect 396579 316644 396580 316708
rect 396644 316644 396645 316708
rect 396579 316643 396645 316644
rect 394739 297396 394805 297397
rect 394739 297332 394740 297396
rect 394804 297332 394805 297396
rect 394739 297331 394805 297332
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 397794 291454 398414 326898
rect 398974 321570 399034 331170
rect 398790 321510 399034 321570
rect 398790 296037 398850 321510
rect 402102 313989 402162 459715
rect 403019 457468 403085 457469
rect 403019 457404 403020 457468
rect 403084 457404 403085 457468
rect 403019 457403 403085 457404
rect 404307 457468 404373 457469
rect 404307 457404 404308 457468
rect 404372 457404 404373 457468
rect 404307 457403 404373 457404
rect 405779 457468 405845 457469
rect 405779 457404 405780 457468
rect 405844 457404 405845 457468
rect 405779 457403 405845 457404
rect 408723 457468 408789 457469
rect 408723 457404 408724 457468
rect 408788 457404 408789 457468
rect 408723 457403 408789 457404
rect 409827 457468 409893 457469
rect 409827 457404 409828 457468
rect 409892 457404 409893 457468
rect 409827 457403 409893 457404
rect 411299 457468 411365 457469
rect 411299 457404 411300 457468
rect 411364 457404 411365 457468
rect 411299 457403 411365 457404
rect 403022 315349 403082 457403
rect 403019 315348 403085 315349
rect 403019 315284 403020 315348
rect 403084 315284 403085 315348
rect 403019 315283 403085 315284
rect 402099 313988 402165 313989
rect 402099 313924 402100 313988
rect 402164 313924 402165 313988
rect 402099 313923 402165 313924
rect 398787 296036 398853 296037
rect 398787 295972 398788 296036
rect 398852 295972 398853 296036
rect 398787 295971 398853 295972
rect 404310 294541 404370 457403
rect 405782 334661 405842 457403
rect 408168 453454 408488 453486
rect 408168 453218 408210 453454
rect 408446 453218 408488 453454
rect 408168 453134 408488 453218
rect 408168 452898 408210 453134
rect 408446 452898 408488 453134
rect 408168 452866 408488 452898
rect 408168 417454 408488 417486
rect 408168 417218 408210 417454
rect 408446 417218 408488 417454
rect 408168 417134 408488 417218
rect 408168 416898 408210 417134
rect 408446 416898 408488 417134
rect 408168 416866 408488 416898
rect 408168 381454 408488 381486
rect 408168 381218 408210 381454
rect 408446 381218 408488 381454
rect 408168 381134 408488 381218
rect 408168 380898 408210 381134
rect 408446 380898 408488 381134
rect 408168 380866 408488 380898
rect 408168 345454 408488 345486
rect 408168 345218 408210 345454
rect 408446 345218 408488 345454
rect 408168 345134 408488 345218
rect 408168 344898 408210 345134
rect 408446 344898 408488 345134
rect 408168 344866 408488 344898
rect 405779 334660 405845 334661
rect 405779 334596 405780 334660
rect 405844 334596 405845 334660
rect 405779 334595 405845 334596
rect 404307 294540 404373 294541
rect 404307 294476 404308 294540
rect 404372 294476 404373 294540
rect 404307 294475 404373 294476
rect 408726 293181 408786 457403
rect 409830 333301 409890 457403
rect 409827 333300 409893 333301
rect 409827 333236 409828 333300
rect 409892 333236 409893 333300
rect 409827 333235 409893 333236
rect 411302 311133 411362 457403
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 411299 311132 411365 311133
rect 411299 311068 411300 311132
rect 411364 311068 411365 311132
rect 411299 311067 411365 311068
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 408723 293180 408789 293181
rect 408723 293116 408724 293180
rect 408788 293116 408789 293180
rect 408723 293115 408789 293116
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 577794 704838 578414 705830
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 254610 453218 254846 453454
rect 254610 452898 254846 453134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 254610 417218 254846 417454
rect 254610 416898 254846 417134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 285330 453218 285566 453454
rect 285330 452898 285566 453134
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 285330 417218 285566 417454
rect 285330 416898 285566 417134
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 316050 453218 316286 453454
rect 316050 452898 316286 453134
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 285330 381218 285566 381454
rect 285330 380898 285566 381134
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 316050 417218 316286 417454
rect 316050 416898 316286 417134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 346770 453218 347006 453454
rect 346770 452898 347006 453134
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 377490 453218 377726 453454
rect 377490 452898 377726 453134
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 361826 435218 362062 435454
rect 362130 435218 362382 435454
rect 361826 434898 362062 435134
rect 362130 434898 362382 435134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 316050 381218 316286 381454
rect 316050 380898 316286 381134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 346770 417218 347006 417454
rect 346770 416898 347006 417134
rect 377490 417218 377726 417454
rect 377490 416898 377726 417134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 361826 399218 362062 399454
rect 362130 399218 362382 399454
rect 361826 398898 362062 399134
rect 362130 398898 362382 399134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 316050 345218 316286 345454
rect 316050 344898 316286 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 346770 381218 347006 381454
rect 346770 380898 347006 381134
rect 377490 381218 377726 381454
rect 377490 380898 377726 381134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 361826 363218 362062 363454
rect 362130 363218 362382 363454
rect 361826 362898 362062 363134
rect 362130 362898 362382 363134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 346770 345218 347006 345454
rect 346770 344898 347006 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 377490 345218 377726 345454
rect 377490 344898 377726 345134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 392850 435218 393086 435454
rect 392850 434898 393086 435134
rect 392850 399218 393086 399454
rect 392850 398898 393086 399134
rect 392850 363218 393086 363454
rect 392850 362898 393086 363134
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 408210 453218 408446 453454
rect 408210 452898 408446 453134
rect 408210 417218 408446 417454
rect 408210 416898 408446 417134
rect 408210 381218 408446 381454
rect 408210 380898 408446 381134
rect 408210 345218 408446 345454
rect 408210 344898 408446 345134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 254610 453454
rect 254846 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 285330 453454
rect 285566 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 316050 453454
rect 316286 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 346770 453454
rect 347006 453218 377490 453454
rect 377726 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 408210 453454
rect 408446 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 254610 453134
rect 254846 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 285330 453134
rect 285566 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 316050 453134
rect 316286 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 346770 453134
rect 347006 452898 377490 453134
rect 377726 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 408210 453134
rect 408446 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 239250 435454
rect 239486 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 269970 435454
rect 270206 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 300690 435454
rect 300926 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 331410 435454
rect 331646 435218 361826 435454
rect 362062 435218 362130 435454
rect 362382 435218 392850 435454
rect 393086 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 239250 435134
rect 239486 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 269970 435134
rect 270206 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 300690 435134
rect 300926 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 331410 435134
rect 331646 434898 361826 435134
rect 362062 434898 362130 435134
rect 362382 434898 392850 435134
rect 393086 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 254610 417454
rect 254846 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 285330 417454
rect 285566 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 316050 417454
rect 316286 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 346770 417454
rect 347006 417218 377490 417454
rect 377726 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 408210 417454
rect 408446 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 254610 417134
rect 254846 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 285330 417134
rect 285566 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 316050 417134
rect 316286 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 346770 417134
rect 347006 416898 377490 417134
rect 377726 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 408210 417134
rect 408446 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 239250 399454
rect 239486 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 269970 399454
rect 270206 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 300690 399454
rect 300926 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 331410 399454
rect 331646 399218 361826 399454
rect 362062 399218 362130 399454
rect 362382 399218 392850 399454
rect 393086 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 239250 399134
rect 239486 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 269970 399134
rect 270206 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 300690 399134
rect 300926 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 331410 399134
rect 331646 398898 361826 399134
rect 362062 398898 362130 399134
rect 362382 398898 392850 399134
rect 393086 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 254610 381454
rect 254846 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 285330 381454
rect 285566 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 316050 381454
rect 316286 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 346770 381454
rect 347006 381218 377490 381454
rect 377726 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 408210 381454
rect 408446 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 254610 381134
rect 254846 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 285330 381134
rect 285566 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 316050 381134
rect 316286 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 346770 381134
rect 347006 380898 377490 381134
rect 377726 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 408210 381134
rect 408446 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 239250 363454
rect 239486 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 269970 363454
rect 270206 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 300690 363454
rect 300926 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 331410 363454
rect 331646 363218 361826 363454
rect 362062 363218 362130 363454
rect 362382 363218 392850 363454
rect 393086 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 239250 363134
rect 239486 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 269970 363134
rect 270206 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 300690 363134
rect 300926 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 331410 363134
rect 331646 362898 361826 363134
rect 362062 362898 362130 363134
rect 362382 362898 392850 363134
rect 393086 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 254610 345454
rect 254846 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 285330 345454
rect 285566 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 316050 345454
rect 316286 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 346770 345454
rect 347006 345218 377490 345454
rect 377726 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 408210 345454
rect 408446 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 254610 345134
rect 254846 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 285330 345134
rect 285566 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 316050 345134
rect 316286 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 346770 345134
rect 347006 344898 377490 345134
rect 377726 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 408210 345134
rect 408446 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use user_proj_example  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box 105 0 179846 120000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 532 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 533 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 535 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 536 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 537 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 538 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 539 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 540 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 541 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 542 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 543 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 544 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 545 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 546 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 547 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 548 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 549 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 550 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 551 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 552 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 553 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 554 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 555 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 556 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 557 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 558 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 559 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 560 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 561 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 562 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 563 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 564 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 565 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 566 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 567 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 568 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 569 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 570 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 571 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 572 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 573 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 574 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 575 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 576 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 577 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 578 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 579 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 580 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 581 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 582 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 583 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 584 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 585 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 586 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 587 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 588 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 589 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 590 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 591 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 592 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 593 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 594 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 595 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 596 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 597 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 598 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 599 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 600 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 601 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 602 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 603 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 604 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 605 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 606 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 607 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 608 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 609 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 610 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 611 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 612 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 613 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 614 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 615 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 616 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 617 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 618 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 619 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 620 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 621 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 622 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 623 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 624 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 625 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 626 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 627 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 628 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 629 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 630 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 631 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 632 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 633 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 634 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 635 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 636 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 637 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
