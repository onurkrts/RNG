magic
tech sky130A
magscale 1 2
timestamp 1647683942
<< obsli1 >>
rect 1104 2159 318872 137649
<< obsm1 >>
rect 290 1096 319594 137680
<< metal2 >>
rect 1398 139200 1454 140000
rect 4158 139200 4214 140000
rect 7010 139200 7066 140000
rect 9770 139200 9826 140000
rect 12622 139200 12678 140000
rect 15382 139200 15438 140000
rect 18234 139200 18290 140000
rect 20994 139200 21050 140000
rect 23846 139200 23902 140000
rect 26606 139200 26662 140000
rect 29458 139200 29514 140000
rect 32218 139200 32274 140000
rect 35070 139200 35126 140000
rect 37830 139200 37886 140000
rect 40682 139200 40738 140000
rect 43442 139200 43498 140000
rect 46294 139200 46350 140000
rect 49054 139200 49110 140000
rect 51906 139200 51962 140000
rect 54666 139200 54722 140000
rect 57518 139200 57574 140000
rect 60278 139200 60334 140000
rect 63130 139200 63186 140000
rect 65890 139200 65946 140000
rect 68742 139200 68798 140000
rect 71502 139200 71558 140000
rect 74354 139200 74410 140000
rect 77114 139200 77170 140000
rect 79966 139200 80022 140000
rect 82726 139200 82782 140000
rect 85578 139200 85634 140000
rect 88338 139200 88394 140000
rect 91190 139200 91246 140000
rect 93950 139200 94006 140000
rect 96802 139200 96858 140000
rect 99562 139200 99618 140000
rect 102414 139200 102470 140000
rect 105174 139200 105230 140000
rect 108026 139200 108082 140000
rect 110786 139200 110842 140000
rect 113638 139200 113694 140000
rect 116398 139200 116454 140000
rect 119250 139200 119306 140000
rect 122010 139200 122066 140000
rect 124862 139200 124918 140000
rect 127622 139200 127678 140000
rect 130474 139200 130530 140000
rect 133234 139200 133290 140000
rect 136086 139200 136142 140000
rect 138846 139200 138902 140000
rect 141698 139200 141754 140000
rect 144458 139200 144514 140000
rect 147310 139200 147366 140000
rect 150070 139200 150126 140000
rect 152922 139200 152978 140000
rect 155682 139200 155738 140000
rect 158534 139200 158590 140000
rect 161386 139200 161442 140000
rect 164146 139200 164202 140000
rect 166998 139200 167054 140000
rect 169758 139200 169814 140000
rect 172610 139200 172666 140000
rect 175370 139200 175426 140000
rect 178222 139200 178278 140000
rect 180982 139200 181038 140000
rect 183834 139200 183890 140000
rect 186594 139200 186650 140000
rect 189446 139200 189502 140000
rect 192206 139200 192262 140000
rect 195058 139200 195114 140000
rect 197818 139200 197874 140000
rect 200670 139200 200726 140000
rect 203430 139200 203486 140000
rect 206282 139200 206338 140000
rect 209042 139200 209098 140000
rect 211894 139200 211950 140000
rect 214654 139200 214710 140000
rect 217506 139200 217562 140000
rect 220266 139200 220322 140000
rect 223118 139200 223174 140000
rect 225878 139200 225934 140000
rect 228730 139200 228786 140000
rect 231490 139200 231546 140000
rect 234342 139200 234398 140000
rect 237102 139200 237158 140000
rect 239954 139200 240010 140000
rect 242714 139200 242770 140000
rect 245566 139200 245622 140000
rect 248326 139200 248382 140000
rect 251178 139200 251234 140000
rect 253938 139200 253994 140000
rect 256790 139200 256846 140000
rect 259550 139200 259606 140000
rect 262402 139200 262458 140000
rect 265162 139200 265218 140000
rect 268014 139200 268070 140000
rect 270774 139200 270830 140000
rect 273626 139200 273682 140000
rect 276386 139200 276442 140000
rect 279238 139200 279294 140000
rect 281998 139200 282054 140000
rect 284850 139200 284906 140000
rect 287610 139200 287666 140000
rect 290462 139200 290518 140000
rect 293222 139200 293278 140000
rect 296074 139200 296130 140000
rect 298834 139200 298890 140000
rect 301686 139200 301742 140000
rect 304446 139200 304502 140000
rect 307298 139200 307354 140000
rect 310058 139200 310114 140000
rect 312910 139200 312966 140000
rect 315670 139200 315726 140000
rect 318522 139200 318578 140000
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2226 0 2282 800
rect 2870 0 2926 800
rect 3514 0 3570 800
rect 4158 0 4214 800
rect 4802 0 4858 800
rect 5446 0 5502 800
rect 6090 0 6146 800
rect 6734 0 6790 800
rect 7378 0 7434 800
rect 8022 0 8078 800
rect 8666 0 8722 800
rect 9310 0 9366 800
rect 9954 0 10010 800
rect 10598 0 10654 800
rect 11242 0 11298 800
rect 11886 0 11942 800
rect 12622 0 12678 800
rect 13266 0 13322 800
rect 13910 0 13966 800
rect 14554 0 14610 800
rect 15198 0 15254 800
rect 15842 0 15898 800
rect 16486 0 16542 800
rect 17130 0 17186 800
rect 17774 0 17830 800
rect 18418 0 18474 800
rect 19062 0 19118 800
rect 19706 0 19762 800
rect 20350 0 20406 800
rect 20994 0 21050 800
rect 21638 0 21694 800
rect 22282 0 22338 800
rect 22926 0 22982 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 24950 0 25006 800
rect 25594 0 25650 800
rect 26238 0 26294 800
rect 26882 0 26938 800
rect 27526 0 27582 800
rect 28170 0 28226 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30102 0 30158 800
rect 30746 0 30802 800
rect 31390 0 31446 800
rect 32034 0 32090 800
rect 32678 0 32734 800
rect 33322 0 33378 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35990 0 36046 800
rect 36634 0 36690 800
rect 37278 0 37334 800
rect 37922 0 37978 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39854 0 39910 800
rect 40498 0 40554 800
rect 41142 0 41198 800
rect 41786 0 41842 800
rect 42430 0 42486 800
rect 43074 0 43130 800
rect 43718 0 43774 800
rect 44362 0 44418 800
rect 45006 0 45062 800
rect 45650 0 45706 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47582 0 47638 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 60002 0 60058 800
rect 60646 0 60702 800
rect 61290 0 61346 800
rect 61934 0 61990 800
rect 62578 0 62634 800
rect 63222 0 63278 800
rect 63866 0 63922 800
rect 64510 0 64566 800
rect 65154 0 65210 800
rect 65798 0 65854 800
rect 66442 0 66498 800
rect 67086 0 67142 800
rect 67730 0 67786 800
rect 68374 0 68430 800
rect 69018 0 69074 800
rect 69662 0 69718 800
rect 70306 0 70362 800
rect 70950 0 71006 800
rect 71686 0 71742 800
rect 72330 0 72386 800
rect 72974 0 73030 800
rect 73618 0 73674 800
rect 74262 0 74318 800
rect 74906 0 74962 800
rect 75550 0 75606 800
rect 76194 0 76250 800
rect 76838 0 76894 800
rect 77482 0 77538 800
rect 78126 0 78182 800
rect 78770 0 78826 800
rect 79414 0 79470 800
rect 80058 0 80114 800
rect 80702 0 80758 800
rect 81346 0 81402 800
rect 81990 0 82046 800
rect 82634 0 82690 800
rect 83370 0 83426 800
rect 84014 0 84070 800
rect 84658 0 84714 800
rect 85302 0 85358 800
rect 85946 0 86002 800
rect 86590 0 86646 800
rect 87234 0 87290 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89166 0 89222 800
rect 89810 0 89866 800
rect 90454 0 90510 800
rect 91098 0 91154 800
rect 91742 0 91798 800
rect 92386 0 92442 800
rect 93030 0 93086 800
rect 93674 0 93730 800
rect 94318 0 94374 800
rect 94962 0 95018 800
rect 95698 0 95754 800
rect 96342 0 96398 800
rect 96986 0 97042 800
rect 97630 0 97686 800
rect 98274 0 98330 800
rect 98918 0 98974 800
rect 99562 0 99618 800
rect 100206 0 100262 800
rect 100850 0 100906 800
rect 101494 0 101550 800
rect 102138 0 102194 800
rect 102782 0 102838 800
rect 103426 0 103482 800
rect 104070 0 104126 800
rect 104714 0 104770 800
rect 105358 0 105414 800
rect 106002 0 106058 800
rect 106646 0 106702 800
rect 107382 0 107438 800
rect 108026 0 108082 800
rect 108670 0 108726 800
rect 109314 0 109370 800
rect 109958 0 110014 800
rect 110602 0 110658 800
rect 111246 0 111302 800
rect 111890 0 111946 800
rect 112534 0 112590 800
rect 113178 0 113234 800
rect 113822 0 113878 800
rect 114466 0 114522 800
rect 115110 0 115166 800
rect 115754 0 115810 800
rect 116398 0 116454 800
rect 117042 0 117098 800
rect 117686 0 117742 800
rect 118330 0 118386 800
rect 119066 0 119122 800
rect 119710 0 119766 800
rect 120354 0 120410 800
rect 120998 0 121054 800
rect 121642 0 121698 800
rect 122286 0 122342 800
rect 122930 0 122986 800
rect 123574 0 123630 800
rect 124218 0 124274 800
rect 124862 0 124918 800
rect 125506 0 125562 800
rect 126150 0 126206 800
rect 126794 0 126850 800
rect 127438 0 127494 800
rect 128082 0 128138 800
rect 128726 0 128782 800
rect 129370 0 129426 800
rect 130014 0 130070 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 133970 0 134026 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139122 0 139178 800
rect 139766 0 139822 800
rect 140410 0 140466 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142342 0 142398 800
rect 143078 0 143134 800
rect 143722 0 143778 800
rect 144366 0 144422 800
rect 145010 0 145066 800
rect 145654 0 145710 800
rect 146298 0 146354 800
rect 146942 0 146998 800
rect 147586 0 147642 800
rect 148230 0 148286 800
rect 148874 0 148930 800
rect 149518 0 149574 800
rect 150162 0 150218 800
rect 150806 0 150862 800
rect 151450 0 151506 800
rect 152094 0 152150 800
rect 152738 0 152794 800
rect 153382 0 153438 800
rect 154026 0 154082 800
rect 154762 0 154818 800
rect 155406 0 155462 800
rect 156050 0 156106 800
rect 156694 0 156750 800
rect 157338 0 157394 800
rect 157982 0 158038 800
rect 158626 0 158682 800
rect 159270 0 159326 800
rect 159914 0 159970 800
rect 160558 0 160614 800
rect 161202 0 161258 800
rect 161846 0 161902 800
rect 162490 0 162546 800
rect 163134 0 163190 800
rect 163778 0 163834 800
rect 164422 0 164478 800
rect 165066 0 165122 800
rect 165710 0 165766 800
rect 166446 0 166502 800
rect 167090 0 167146 800
rect 167734 0 167790 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169666 0 169722 800
rect 170310 0 170366 800
rect 170954 0 171010 800
rect 171598 0 171654 800
rect 172242 0 172298 800
rect 172886 0 172942 800
rect 173530 0 173586 800
rect 174174 0 174230 800
rect 174818 0 174874 800
rect 175462 0 175518 800
rect 176106 0 176162 800
rect 176750 0 176806 800
rect 177394 0 177450 800
rect 178130 0 178186 800
rect 178774 0 178830 800
rect 179418 0 179474 800
rect 180062 0 180118 800
rect 180706 0 180762 800
rect 181350 0 181406 800
rect 181994 0 182050 800
rect 182638 0 182694 800
rect 183282 0 183338 800
rect 183926 0 183982 800
rect 184570 0 184626 800
rect 185214 0 185270 800
rect 185858 0 185914 800
rect 186502 0 186558 800
rect 187146 0 187202 800
rect 187790 0 187846 800
rect 188434 0 188490 800
rect 189078 0 189134 800
rect 189722 0 189778 800
rect 190458 0 190514 800
rect 191102 0 191158 800
rect 191746 0 191802 800
rect 192390 0 192446 800
rect 193034 0 193090 800
rect 193678 0 193734 800
rect 194322 0 194378 800
rect 194966 0 195022 800
rect 195610 0 195666 800
rect 196254 0 196310 800
rect 196898 0 196954 800
rect 197542 0 197598 800
rect 198186 0 198242 800
rect 198830 0 198886 800
rect 199474 0 199530 800
rect 200118 0 200174 800
rect 200762 0 200818 800
rect 201406 0 201462 800
rect 202142 0 202198 800
rect 202786 0 202842 800
rect 203430 0 203486 800
rect 204074 0 204130 800
rect 204718 0 204774 800
rect 205362 0 205418 800
rect 206006 0 206062 800
rect 206650 0 206706 800
rect 207294 0 207350 800
rect 207938 0 207994 800
rect 208582 0 208638 800
rect 209226 0 209282 800
rect 209870 0 209926 800
rect 210514 0 210570 800
rect 211158 0 211214 800
rect 211802 0 211858 800
rect 212446 0 212502 800
rect 213090 0 213146 800
rect 213826 0 213882 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215758 0 215814 800
rect 216402 0 216458 800
rect 217046 0 217102 800
rect 217690 0 217746 800
rect 218334 0 218390 800
rect 218978 0 219034 800
rect 219622 0 219678 800
rect 220266 0 220322 800
rect 220910 0 220966 800
rect 221554 0 221610 800
rect 222198 0 222254 800
rect 222842 0 222898 800
rect 223486 0 223542 800
rect 224130 0 224186 800
rect 224774 0 224830 800
rect 225510 0 225566 800
rect 226154 0 226210 800
rect 226798 0 226854 800
rect 227442 0 227498 800
rect 228086 0 228142 800
rect 228730 0 228786 800
rect 229374 0 229430 800
rect 230018 0 230074 800
rect 230662 0 230718 800
rect 231306 0 231362 800
rect 231950 0 232006 800
rect 232594 0 232650 800
rect 233238 0 233294 800
rect 233882 0 233938 800
rect 234526 0 234582 800
rect 235170 0 235226 800
rect 235814 0 235870 800
rect 236458 0 236514 800
rect 237102 0 237158 800
rect 237838 0 237894 800
rect 238482 0 238538 800
rect 239126 0 239182 800
rect 239770 0 239826 800
rect 240414 0 240470 800
rect 241058 0 241114 800
rect 241702 0 241758 800
rect 242346 0 242402 800
rect 242990 0 243046 800
rect 243634 0 243690 800
rect 244278 0 244334 800
rect 244922 0 244978 800
rect 245566 0 245622 800
rect 246210 0 246266 800
rect 246854 0 246910 800
rect 247498 0 247554 800
rect 248142 0 248198 800
rect 248786 0 248842 800
rect 249522 0 249578 800
rect 250166 0 250222 800
rect 250810 0 250866 800
rect 251454 0 251510 800
rect 252098 0 252154 800
rect 252742 0 252798 800
rect 253386 0 253442 800
rect 254030 0 254086 800
rect 254674 0 254730 800
rect 255318 0 255374 800
rect 255962 0 256018 800
rect 256606 0 256662 800
rect 257250 0 257306 800
rect 257894 0 257950 800
rect 258538 0 258594 800
rect 259182 0 259238 800
rect 259826 0 259882 800
rect 260470 0 260526 800
rect 261206 0 261262 800
rect 261850 0 261906 800
rect 262494 0 262550 800
rect 263138 0 263194 800
rect 263782 0 263838 800
rect 264426 0 264482 800
rect 265070 0 265126 800
rect 265714 0 265770 800
rect 266358 0 266414 800
rect 267002 0 267058 800
rect 267646 0 267702 800
rect 268290 0 268346 800
rect 268934 0 268990 800
rect 269578 0 269634 800
rect 270222 0 270278 800
rect 270866 0 270922 800
rect 271510 0 271566 800
rect 272154 0 272210 800
rect 272890 0 272946 800
rect 273534 0 273590 800
rect 274178 0 274234 800
rect 274822 0 274878 800
rect 275466 0 275522 800
rect 276110 0 276166 800
rect 276754 0 276810 800
rect 277398 0 277454 800
rect 278042 0 278098 800
rect 278686 0 278742 800
rect 279330 0 279386 800
rect 279974 0 280030 800
rect 280618 0 280674 800
rect 281262 0 281318 800
rect 281906 0 281962 800
rect 282550 0 282606 800
rect 283194 0 283250 800
rect 283838 0 283894 800
rect 284482 0 284538 800
rect 285218 0 285274 800
rect 285862 0 285918 800
rect 286506 0 286562 800
rect 287150 0 287206 800
rect 287794 0 287850 800
rect 288438 0 288494 800
rect 289082 0 289138 800
rect 289726 0 289782 800
rect 290370 0 290426 800
rect 291014 0 291070 800
rect 291658 0 291714 800
rect 292302 0 292358 800
rect 292946 0 293002 800
rect 293590 0 293646 800
rect 294234 0 294290 800
rect 294878 0 294934 800
rect 295522 0 295578 800
rect 296166 0 296222 800
rect 296902 0 296958 800
rect 297546 0 297602 800
rect 298190 0 298246 800
rect 298834 0 298890 800
rect 299478 0 299534 800
rect 300122 0 300178 800
rect 300766 0 300822 800
rect 301410 0 301466 800
rect 302054 0 302110 800
rect 302698 0 302754 800
rect 303342 0 303398 800
rect 303986 0 304042 800
rect 304630 0 304686 800
rect 305274 0 305330 800
rect 305918 0 305974 800
rect 306562 0 306618 800
rect 307206 0 307262 800
rect 307850 0 307906 800
rect 308586 0 308642 800
rect 309230 0 309286 800
rect 309874 0 309930 800
rect 310518 0 310574 800
rect 311162 0 311218 800
rect 311806 0 311862 800
rect 312450 0 312506 800
rect 313094 0 313150 800
rect 313738 0 313794 800
rect 314382 0 314438 800
rect 315026 0 315082 800
rect 315670 0 315726 800
rect 316314 0 316370 800
rect 316958 0 317014 800
rect 317602 0 317658 800
rect 318246 0 318302 800
rect 318890 0 318946 800
rect 319534 0 319590 800
<< obsm2 >>
rect 296 139144 1342 139346
rect 1510 139144 4102 139346
rect 4270 139144 6954 139346
rect 7122 139144 9714 139346
rect 9882 139144 12566 139346
rect 12734 139144 15326 139346
rect 15494 139144 18178 139346
rect 18346 139144 20938 139346
rect 21106 139144 23790 139346
rect 23958 139144 26550 139346
rect 26718 139144 29402 139346
rect 29570 139144 32162 139346
rect 32330 139144 35014 139346
rect 35182 139144 37774 139346
rect 37942 139144 40626 139346
rect 40794 139144 43386 139346
rect 43554 139144 46238 139346
rect 46406 139144 48998 139346
rect 49166 139144 51850 139346
rect 52018 139144 54610 139346
rect 54778 139144 57462 139346
rect 57630 139144 60222 139346
rect 60390 139144 63074 139346
rect 63242 139144 65834 139346
rect 66002 139144 68686 139346
rect 68854 139144 71446 139346
rect 71614 139144 74298 139346
rect 74466 139144 77058 139346
rect 77226 139144 79910 139346
rect 80078 139144 82670 139346
rect 82838 139144 85522 139346
rect 85690 139144 88282 139346
rect 88450 139144 91134 139346
rect 91302 139144 93894 139346
rect 94062 139144 96746 139346
rect 96914 139144 99506 139346
rect 99674 139144 102358 139346
rect 102526 139144 105118 139346
rect 105286 139144 107970 139346
rect 108138 139144 110730 139346
rect 110898 139144 113582 139346
rect 113750 139144 116342 139346
rect 116510 139144 119194 139346
rect 119362 139144 121954 139346
rect 122122 139144 124806 139346
rect 124974 139144 127566 139346
rect 127734 139144 130418 139346
rect 130586 139144 133178 139346
rect 133346 139144 136030 139346
rect 136198 139144 138790 139346
rect 138958 139144 141642 139346
rect 141810 139144 144402 139346
rect 144570 139144 147254 139346
rect 147422 139144 150014 139346
rect 150182 139144 152866 139346
rect 153034 139144 155626 139346
rect 155794 139144 158478 139346
rect 158646 139144 161330 139346
rect 161498 139144 164090 139346
rect 164258 139144 166942 139346
rect 167110 139144 169702 139346
rect 169870 139144 172554 139346
rect 172722 139144 175314 139346
rect 175482 139144 178166 139346
rect 178334 139144 180926 139346
rect 181094 139144 183778 139346
rect 183946 139144 186538 139346
rect 186706 139144 189390 139346
rect 189558 139144 192150 139346
rect 192318 139144 195002 139346
rect 195170 139144 197762 139346
rect 197930 139144 200614 139346
rect 200782 139144 203374 139346
rect 203542 139144 206226 139346
rect 206394 139144 208986 139346
rect 209154 139144 211838 139346
rect 212006 139144 214598 139346
rect 214766 139144 217450 139346
rect 217618 139144 220210 139346
rect 220378 139144 223062 139346
rect 223230 139144 225822 139346
rect 225990 139144 228674 139346
rect 228842 139144 231434 139346
rect 231602 139144 234286 139346
rect 234454 139144 237046 139346
rect 237214 139144 239898 139346
rect 240066 139144 242658 139346
rect 242826 139144 245510 139346
rect 245678 139144 248270 139346
rect 248438 139144 251122 139346
rect 251290 139144 253882 139346
rect 254050 139144 256734 139346
rect 256902 139144 259494 139346
rect 259662 139144 262346 139346
rect 262514 139144 265106 139346
rect 265274 139144 267958 139346
rect 268126 139144 270718 139346
rect 270886 139144 273570 139346
rect 273738 139144 276330 139346
rect 276498 139144 279182 139346
rect 279350 139144 281942 139346
rect 282110 139144 284794 139346
rect 284962 139144 287554 139346
rect 287722 139144 290406 139346
rect 290574 139144 293166 139346
rect 293334 139144 296018 139346
rect 296186 139144 298778 139346
rect 298946 139144 301630 139346
rect 301798 139144 304390 139346
rect 304558 139144 307242 139346
rect 307410 139144 310002 139346
rect 310170 139144 312854 139346
rect 313022 139144 315614 139346
rect 315782 139144 318466 139346
rect 318634 139144 319588 139346
rect 296 856 319588 139144
rect 406 734 882 856
rect 1050 734 1526 856
rect 1694 734 2170 856
rect 2338 734 2814 856
rect 2982 734 3458 856
rect 3626 734 4102 856
rect 4270 734 4746 856
rect 4914 734 5390 856
rect 5558 734 6034 856
rect 6202 734 6678 856
rect 6846 734 7322 856
rect 7490 734 7966 856
rect 8134 734 8610 856
rect 8778 734 9254 856
rect 9422 734 9898 856
rect 10066 734 10542 856
rect 10710 734 11186 856
rect 11354 734 11830 856
rect 11998 734 12566 856
rect 12734 734 13210 856
rect 13378 734 13854 856
rect 14022 734 14498 856
rect 14666 734 15142 856
rect 15310 734 15786 856
rect 15954 734 16430 856
rect 16598 734 17074 856
rect 17242 734 17718 856
rect 17886 734 18362 856
rect 18530 734 19006 856
rect 19174 734 19650 856
rect 19818 734 20294 856
rect 20462 734 20938 856
rect 21106 734 21582 856
rect 21750 734 22226 856
rect 22394 734 22870 856
rect 23038 734 23514 856
rect 23682 734 24250 856
rect 24418 734 24894 856
rect 25062 734 25538 856
rect 25706 734 26182 856
rect 26350 734 26826 856
rect 26994 734 27470 856
rect 27638 734 28114 856
rect 28282 734 28758 856
rect 28926 734 29402 856
rect 29570 734 30046 856
rect 30214 734 30690 856
rect 30858 734 31334 856
rect 31502 734 31978 856
rect 32146 734 32622 856
rect 32790 734 33266 856
rect 33434 734 33910 856
rect 34078 734 34554 856
rect 34722 734 35198 856
rect 35366 734 35934 856
rect 36102 734 36578 856
rect 36746 734 37222 856
rect 37390 734 37866 856
rect 38034 734 38510 856
rect 38678 734 39154 856
rect 39322 734 39798 856
rect 39966 734 40442 856
rect 40610 734 41086 856
rect 41254 734 41730 856
rect 41898 734 42374 856
rect 42542 734 43018 856
rect 43186 734 43662 856
rect 43830 734 44306 856
rect 44474 734 44950 856
rect 45118 734 45594 856
rect 45762 734 46238 856
rect 46406 734 46882 856
rect 47050 734 47526 856
rect 47694 734 48262 856
rect 48430 734 48906 856
rect 49074 734 49550 856
rect 49718 734 50194 856
rect 50362 734 50838 856
rect 51006 734 51482 856
rect 51650 734 52126 856
rect 52294 734 52770 856
rect 52938 734 53414 856
rect 53582 734 54058 856
rect 54226 734 54702 856
rect 54870 734 55346 856
rect 55514 734 55990 856
rect 56158 734 56634 856
rect 56802 734 57278 856
rect 57446 734 57922 856
rect 58090 734 58566 856
rect 58734 734 59210 856
rect 59378 734 59946 856
rect 60114 734 60590 856
rect 60758 734 61234 856
rect 61402 734 61878 856
rect 62046 734 62522 856
rect 62690 734 63166 856
rect 63334 734 63810 856
rect 63978 734 64454 856
rect 64622 734 65098 856
rect 65266 734 65742 856
rect 65910 734 66386 856
rect 66554 734 67030 856
rect 67198 734 67674 856
rect 67842 734 68318 856
rect 68486 734 68962 856
rect 69130 734 69606 856
rect 69774 734 70250 856
rect 70418 734 70894 856
rect 71062 734 71630 856
rect 71798 734 72274 856
rect 72442 734 72918 856
rect 73086 734 73562 856
rect 73730 734 74206 856
rect 74374 734 74850 856
rect 75018 734 75494 856
rect 75662 734 76138 856
rect 76306 734 76782 856
rect 76950 734 77426 856
rect 77594 734 78070 856
rect 78238 734 78714 856
rect 78882 734 79358 856
rect 79526 734 80002 856
rect 80170 734 80646 856
rect 80814 734 81290 856
rect 81458 734 81934 856
rect 82102 734 82578 856
rect 82746 734 83314 856
rect 83482 734 83958 856
rect 84126 734 84602 856
rect 84770 734 85246 856
rect 85414 734 85890 856
rect 86058 734 86534 856
rect 86702 734 87178 856
rect 87346 734 87822 856
rect 87990 734 88466 856
rect 88634 734 89110 856
rect 89278 734 89754 856
rect 89922 734 90398 856
rect 90566 734 91042 856
rect 91210 734 91686 856
rect 91854 734 92330 856
rect 92498 734 92974 856
rect 93142 734 93618 856
rect 93786 734 94262 856
rect 94430 734 94906 856
rect 95074 734 95642 856
rect 95810 734 96286 856
rect 96454 734 96930 856
rect 97098 734 97574 856
rect 97742 734 98218 856
rect 98386 734 98862 856
rect 99030 734 99506 856
rect 99674 734 100150 856
rect 100318 734 100794 856
rect 100962 734 101438 856
rect 101606 734 102082 856
rect 102250 734 102726 856
rect 102894 734 103370 856
rect 103538 734 104014 856
rect 104182 734 104658 856
rect 104826 734 105302 856
rect 105470 734 105946 856
rect 106114 734 106590 856
rect 106758 734 107326 856
rect 107494 734 107970 856
rect 108138 734 108614 856
rect 108782 734 109258 856
rect 109426 734 109902 856
rect 110070 734 110546 856
rect 110714 734 111190 856
rect 111358 734 111834 856
rect 112002 734 112478 856
rect 112646 734 113122 856
rect 113290 734 113766 856
rect 113934 734 114410 856
rect 114578 734 115054 856
rect 115222 734 115698 856
rect 115866 734 116342 856
rect 116510 734 116986 856
rect 117154 734 117630 856
rect 117798 734 118274 856
rect 118442 734 119010 856
rect 119178 734 119654 856
rect 119822 734 120298 856
rect 120466 734 120942 856
rect 121110 734 121586 856
rect 121754 734 122230 856
rect 122398 734 122874 856
rect 123042 734 123518 856
rect 123686 734 124162 856
rect 124330 734 124806 856
rect 124974 734 125450 856
rect 125618 734 126094 856
rect 126262 734 126738 856
rect 126906 734 127382 856
rect 127550 734 128026 856
rect 128194 734 128670 856
rect 128838 734 129314 856
rect 129482 734 129958 856
rect 130126 734 130694 856
rect 130862 734 131338 856
rect 131506 734 131982 856
rect 132150 734 132626 856
rect 132794 734 133270 856
rect 133438 734 133914 856
rect 134082 734 134558 856
rect 134726 734 135202 856
rect 135370 734 135846 856
rect 136014 734 136490 856
rect 136658 734 137134 856
rect 137302 734 137778 856
rect 137946 734 138422 856
rect 138590 734 139066 856
rect 139234 734 139710 856
rect 139878 734 140354 856
rect 140522 734 140998 856
rect 141166 734 141642 856
rect 141810 734 142286 856
rect 142454 734 143022 856
rect 143190 734 143666 856
rect 143834 734 144310 856
rect 144478 734 144954 856
rect 145122 734 145598 856
rect 145766 734 146242 856
rect 146410 734 146886 856
rect 147054 734 147530 856
rect 147698 734 148174 856
rect 148342 734 148818 856
rect 148986 734 149462 856
rect 149630 734 150106 856
rect 150274 734 150750 856
rect 150918 734 151394 856
rect 151562 734 152038 856
rect 152206 734 152682 856
rect 152850 734 153326 856
rect 153494 734 153970 856
rect 154138 734 154706 856
rect 154874 734 155350 856
rect 155518 734 155994 856
rect 156162 734 156638 856
rect 156806 734 157282 856
rect 157450 734 157926 856
rect 158094 734 158570 856
rect 158738 734 159214 856
rect 159382 734 159858 856
rect 160026 734 160502 856
rect 160670 734 161146 856
rect 161314 734 161790 856
rect 161958 734 162434 856
rect 162602 734 163078 856
rect 163246 734 163722 856
rect 163890 734 164366 856
rect 164534 734 165010 856
rect 165178 734 165654 856
rect 165822 734 166390 856
rect 166558 734 167034 856
rect 167202 734 167678 856
rect 167846 734 168322 856
rect 168490 734 168966 856
rect 169134 734 169610 856
rect 169778 734 170254 856
rect 170422 734 170898 856
rect 171066 734 171542 856
rect 171710 734 172186 856
rect 172354 734 172830 856
rect 172998 734 173474 856
rect 173642 734 174118 856
rect 174286 734 174762 856
rect 174930 734 175406 856
rect 175574 734 176050 856
rect 176218 734 176694 856
rect 176862 734 177338 856
rect 177506 734 178074 856
rect 178242 734 178718 856
rect 178886 734 179362 856
rect 179530 734 180006 856
rect 180174 734 180650 856
rect 180818 734 181294 856
rect 181462 734 181938 856
rect 182106 734 182582 856
rect 182750 734 183226 856
rect 183394 734 183870 856
rect 184038 734 184514 856
rect 184682 734 185158 856
rect 185326 734 185802 856
rect 185970 734 186446 856
rect 186614 734 187090 856
rect 187258 734 187734 856
rect 187902 734 188378 856
rect 188546 734 189022 856
rect 189190 734 189666 856
rect 189834 734 190402 856
rect 190570 734 191046 856
rect 191214 734 191690 856
rect 191858 734 192334 856
rect 192502 734 192978 856
rect 193146 734 193622 856
rect 193790 734 194266 856
rect 194434 734 194910 856
rect 195078 734 195554 856
rect 195722 734 196198 856
rect 196366 734 196842 856
rect 197010 734 197486 856
rect 197654 734 198130 856
rect 198298 734 198774 856
rect 198942 734 199418 856
rect 199586 734 200062 856
rect 200230 734 200706 856
rect 200874 734 201350 856
rect 201518 734 202086 856
rect 202254 734 202730 856
rect 202898 734 203374 856
rect 203542 734 204018 856
rect 204186 734 204662 856
rect 204830 734 205306 856
rect 205474 734 205950 856
rect 206118 734 206594 856
rect 206762 734 207238 856
rect 207406 734 207882 856
rect 208050 734 208526 856
rect 208694 734 209170 856
rect 209338 734 209814 856
rect 209982 734 210458 856
rect 210626 734 211102 856
rect 211270 734 211746 856
rect 211914 734 212390 856
rect 212558 734 213034 856
rect 213202 734 213770 856
rect 213938 734 214414 856
rect 214582 734 215058 856
rect 215226 734 215702 856
rect 215870 734 216346 856
rect 216514 734 216990 856
rect 217158 734 217634 856
rect 217802 734 218278 856
rect 218446 734 218922 856
rect 219090 734 219566 856
rect 219734 734 220210 856
rect 220378 734 220854 856
rect 221022 734 221498 856
rect 221666 734 222142 856
rect 222310 734 222786 856
rect 222954 734 223430 856
rect 223598 734 224074 856
rect 224242 734 224718 856
rect 224886 734 225454 856
rect 225622 734 226098 856
rect 226266 734 226742 856
rect 226910 734 227386 856
rect 227554 734 228030 856
rect 228198 734 228674 856
rect 228842 734 229318 856
rect 229486 734 229962 856
rect 230130 734 230606 856
rect 230774 734 231250 856
rect 231418 734 231894 856
rect 232062 734 232538 856
rect 232706 734 233182 856
rect 233350 734 233826 856
rect 233994 734 234470 856
rect 234638 734 235114 856
rect 235282 734 235758 856
rect 235926 734 236402 856
rect 236570 734 237046 856
rect 237214 734 237782 856
rect 237950 734 238426 856
rect 238594 734 239070 856
rect 239238 734 239714 856
rect 239882 734 240358 856
rect 240526 734 241002 856
rect 241170 734 241646 856
rect 241814 734 242290 856
rect 242458 734 242934 856
rect 243102 734 243578 856
rect 243746 734 244222 856
rect 244390 734 244866 856
rect 245034 734 245510 856
rect 245678 734 246154 856
rect 246322 734 246798 856
rect 246966 734 247442 856
rect 247610 734 248086 856
rect 248254 734 248730 856
rect 248898 734 249466 856
rect 249634 734 250110 856
rect 250278 734 250754 856
rect 250922 734 251398 856
rect 251566 734 252042 856
rect 252210 734 252686 856
rect 252854 734 253330 856
rect 253498 734 253974 856
rect 254142 734 254618 856
rect 254786 734 255262 856
rect 255430 734 255906 856
rect 256074 734 256550 856
rect 256718 734 257194 856
rect 257362 734 257838 856
rect 258006 734 258482 856
rect 258650 734 259126 856
rect 259294 734 259770 856
rect 259938 734 260414 856
rect 260582 734 261150 856
rect 261318 734 261794 856
rect 261962 734 262438 856
rect 262606 734 263082 856
rect 263250 734 263726 856
rect 263894 734 264370 856
rect 264538 734 265014 856
rect 265182 734 265658 856
rect 265826 734 266302 856
rect 266470 734 266946 856
rect 267114 734 267590 856
rect 267758 734 268234 856
rect 268402 734 268878 856
rect 269046 734 269522 856
rect 269690 734 270166 856
rect 270334 734 270810 856
rect 270978 734 271454 856
rect 271622 734 272098 856
rect 272266 734 272834 856
rect 273002 734 273478 856
rect 273646 734 274122 856
rect 274290 734 274766 856
rect 274934 734 275410 856
rect 275578 734 276054 856
rect 276222 734 276698 856
rect 276866 734 277342 856
rect 277510 734 277986 856
rect 278154 734 278630 856
rect 278798 734 279274 856
rect 279442 734 279918 856
rect 280086 734 280562 856
rect 280730 734 281206 856
rect 281374 734 281850 856
rect 282018 734 282494 856
rect 282662 734 283138 856
rect 283306 734 283782 856
rect 283950 734 284426 856
rect 284594 734 285162 856
rect 285330 734 285806 856
rect 285974 734 286450 856
rect 286618 734 287094 856
rect 287262 734 287738 856
rect 287906 734 288382 856
rect 288550 734 289026 856
rect 289194 734 289670 856
rect 289838 734 290314 856
rect 290482 734 290958 856
rect 291126 734 291602 856
rect 291770 734 292246 856
rect 292414 734 292890 856
rect 293058 734 293534 856
rect 293702 734 294178 856
rect 294346 734 294822 856
rect 294990 734 295466 856
rect 295634 734 296110 856
rect 296278 734 296846 856
rect 297014 734 297490 856
rect 297658 734 298134 856
rect 298302 734 298778 856
rect 298946 734 299422 856
rect 299590 734 300066 856
rect 300234 734 300710 856
rect 300878 734 301354 856
rect 301522 734 301998 856
rect 302166 734 302642 856
rect 302810 734 303286 856
rect 303454 734 303930 856
rect 304098 734 304574 856
rect 304742 734 305218 856
rect 305386 734 305862 856
rect 306030 734 306506 856
rect 306674 734 307150 856
rect 307318 734 307794 856
rect 307962 734 308530 856
rect 308698 734 309174 856
rect 309342 734 309818 856
rect 309986 734 310462 856
rect 310630 734 311106 856
rect 311274 734 311750 856
rect 311918 734 312394 856
rect 312562 734 313038 856
rect 313206 734 313682 856
rect 313850 734 314326 856
rect 314494 734 314970 856
rect 315138 734 315614 856
rect 315782 734 316258 856
rect 316426 734 316902 856
rect 317070 734 317546 856
rect 317714 734 318190 856
rect 318358 734 318834 856
rect 319002 734 319478 856
<< obsm3 >>
rect 4208 1259 314528 137665
<< metal4 >>
rect 4208 2128 4528 137680
rect 14208 2128 14528 137680
rect 24208 2128 24528 137680
rect 34208 2128 34528 137680
rect 44208 2128 44528 137680
rect 54208 2128 54528 137680
rect 64208 2128 64528 137680
rect 74208 2128 74528 137680
rect 84208 2128 84528 137680
rect 94208 2128 94528 137680
rect 104208 2128 104528 137680
rect 114208 2128 114528 137680
rect 124208 2128 124528 137680
rect 134208 2128 134528 137680
rect 144208 2128 144528 137680
rect 154208 2128 154528 137680
rect 164208 2128 164528 137680
rect 174208 2128 174528 137680
rect 184208 2128 184528 137680
rect 194208 2128 194528 137680
rect 204208 2128 204528 137680
rect 214208 2128 214528 137680
rect 224208 2128 224528 137680
rect 234208 2128 234528 137680
rect 244208 2128 244528 137680
rect 254208 2128 254528 137680
rect 264208 2128 264528 137680
rect 274208 2128 274528 137680
rect 284208 2128 284528 137680
rect 294208 2128 294528 137680
rect 304208 2128 304528 137680
rect 314208 2128 314528 137680
<< obsm4 >>
rect 144683 3163 154128 14381
rect 154608 3163 164128 14381
rect 164608 3163 174128 14381
rect 174608 3163 184128 14381
rect 184608 3163 192405 14381
<< labels >>
rlabel metal2 s 1398 139200 1454 140000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 85578 139200 85634 140000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 93950 139200 94006 140000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 102414 139200 102470 140000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 110786 139200 110842 140000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 119250 139200 119306 140000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 127622 139200 127678 140000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 136086 139200 136142 140000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 144458 139200 144514 140000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 152922 139200 152978 140000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 161386 139200 161442 140000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 9770 139200 9826 140000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 169758 139200 169814 140000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 178222 139200 178278 140000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 186594 139200 186650 140000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 195058 139200 195114 140000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 203430 139200 203486 140000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 211894 139200 211950 140000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 220266 139200 220322 140000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 228730 139200 228786 140000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 237102 139200 237158 140000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 245566 139200 245622 140000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 18234 139200 18290 140000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 253938 139200 253994 140000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 262402 139200 262458 140000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 270774 139200 270830 140000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 279238 139200 279294 140000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 287610 139200 287666 140000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 296074 139200 296130 140000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 304446 139200 304502 140000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 312910 139200 312966 140000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 26606 139200 26662 140000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 35070 139200 35126 140000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 43442 139200 43498 140000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 51906 139200 51962 140000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 60278 139200 60334 140000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 68742 139200 68798 140000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 77114 139200 77170 140000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4158 139200 4214 140000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 88338 139200 88394 140000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 96802 139200 96858 140000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 105174 139200 105230 140000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 113638 139200 113694 140000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 122010 139200 122066 140000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 130474 139200 130530 140000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 138846 139200 138902 140000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 147310 139200 147366 140000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 155682 139200 155738 140000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 164146 139200 164202 140000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 12622 139200 12678 140000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 172610 139200 172666 140000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 180982 139200 181038 140000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 189446 139200 189502 140000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 197818 139200 197874 140000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 206282 139200 206338 140000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 214654 139200 214710 140000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 223118 139200 223174 140000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 231490 139200 231546 140000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 239954 139200 240010 140000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 248326 139200 248382 140000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 20994 139200 21050 140000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 256790 139200 256846 140000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 265162 139200 265218 140000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 273626 139200 273682 140000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 281998 139200 282054 140000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 290462 139200 290518 140000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 298834 139200 298890 140000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 307298 139200 307354 140000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 315670 139200 315726 140000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 29458 139200 29514 140000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 37830 139200 37886 140000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 46294 139200 46350 140000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 54666 139200 54722 140000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 63130 139200 63186 140000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 71502 139200 71558 140000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 79966 139200 80022 140000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 7010 139200 7066 140000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 91190 139200 91246 140000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 99562 139200 99618 140000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 108026 139200 108082 140000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 116398 139200 116454 140000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 124862 139200 124918 140000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 133234 139200 133290 140000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 141698 139200 141754 140000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 150070 139200 150126 140000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 158534 139200 158590 140000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 166998 139200 167054 140000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 15382 139200 15438 140000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 175370 139200 175426 140000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 183834 139200 183890 140000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 192206 139200 192262 140000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 200670 139200 200726 140000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 209042 139200 209098 140000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 217506 139200 217562 140000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 225878 139200 225934 140000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 234342 139200 234398 140000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 242714 139200 242770 140000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 251178 139200 251234 140000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 23846 139200 23902 140000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 259550 139200 259606 140000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 268014 139200 268070 140000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 276386 139200 276442 140000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 284850 139200 284906 140000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 293222 139200 293278 140000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 301686 139200 301742 140000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 310058 139200 310114 140000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 318522 139200 318578 140000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 32218 139200 32274 140000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 40682 139200 40738 140000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 49054 139200 49110 140000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 57518 139200 57574 140000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 65890 139200 65946 140000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 74354 139200 74410 140000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 82726 139200 82782 140000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 318246 0 318302 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 318890 0 318946 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 319534 0 319590 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 265714 0 265770 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 267646 0 267702 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 269578 0 269634 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 271510 0 271566 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 273534 0 273590 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 277398 0 277454 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 279330 0 279386 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 281262 0 281318 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 283194 0 283250 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 287150 0 287206 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 292946 0 293002 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 298834 0 298890 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 306562 0 306618 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 308586 0 308642 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 310518 0 310574 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 312450 0 312506 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 316314 0 316370 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 181994 0 182050 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 199474 0 199530 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 201406 0 201462 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 207294 0 207350 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 209226 0 209282 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 211158 0 211214 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 213090 0 213146 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 228730 0 228786 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 232594 0 232650 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 238482 0 238538 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 242346 0 242402 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 246210 0 246266 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 259826 0 259882 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 264426 0 264482 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 266358 0 266414 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 268290 0 268346 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 270222 0 270278 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 272154 0 272210 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 274178 0 274234 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 276110 0 276166 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 278042 0 278098 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 279974 0 280030 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 283838 0 283894 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 285862 0 285918 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 287794 0 287850 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 289726 0 289782 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 291658 0 291714 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 293590 0 293646 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 295522 0 295578 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 297546 0 297602 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 299478 0 299534 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 301410 0 301466 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 303342 0 303398 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 305274 0 305330 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 307206 0 307262 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 309230 0 309286 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 313094 0 313150 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 315026 0 315082 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 316958 0 317014 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 170954 0 171010 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 178774 0 178830 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 182638 0 182694 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 186502 0 186558 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 190458 0 190514 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 192390 0 192446 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 196254 0 196310 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 198186 0 198242 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 200118 0 200174 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 202142 0 202198 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 206006 0 206062 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 207938 0 207994 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 209870 0 209926 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 211802 0 211858 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 215758 0 215814 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 225510 0 225566 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 227442 0 227498 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 229374 0 229430 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 231306 0 231362 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 233238 0 233294 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 235170 0 235226 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 237102 0 237158 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 239126 0 239182 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 244922 0 244978 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 246854 0 246910 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 248786 0 248842 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 250810 0 250866 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 258538 0 258594 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 262494 0 262550 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 265070 0 265126 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 270866 0 270922 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 274822 0 274878 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 278686 0 278742 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 282550 0 282606 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 284482 0 284538 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 286506 0 286562 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 288438 0 288494 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 292302 0 292358 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 294234 0 294290 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 296166 0 296222 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 302054 0 302110 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 303986 0 304042 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 305918 0 305974 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 309874 0 309930 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 313738 0 313794 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 315670 0 315726 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 198830 0 198886 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 220266 0 220322 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 226154 0 226210 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 231950 0 232006 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 255318 0 255374 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 261206 0 261262 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 24208 2128 24528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 44208 2128 44528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 64208 2128 64528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 84208 2128 84528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 104208 2128 104528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 124208 2128 124528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 144208 2128 144528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 164208 2128 164528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 184208 2128 184528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 204208 2128 204528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 224208 2128 224528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 244208 2128 244528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 264208 2128 264528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 284208 2128 284528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 304208 2128 304528 137680 6 vccd1
port 502 nsew power input
rlabel metal4 s 14208 2128 14528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 34208 2128 34528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 54208 2128 54528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 74208 2128 74528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 94208 2128 94528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 114208 2128 114528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 134208 2128 134528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 154208 2128 154528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 174208 2128 174528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 194208 2128 194528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 214208 2128 214528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234208 2128 234528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 254208 2128 254528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 274208 2128 274528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 294208 2128 294528 137680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 314208 2128 314528 137680 6 vssd1
port 503 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 320000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18400186
string GDS_FILE /home/asrock/caravel_tutorial/RNG/openlane/rng_chaos/runs/rng_chaos/results/finishing/rng_chaos_top.magic.gds
string GDS_START 794350
<< end >>

