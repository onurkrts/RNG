magic
tech sky130A
magscale 1 2
timestamp 1647848066
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 283834 700816 283840 700868
rect 283892 700856 283898 700868
rect 328454 700856 328460 700868
rect 283892 700828 328460 700856
rect 283892 700816 283898 700828
rect 328454 700816 328460 700828
rect 328512 700816 328518 700868
rect 318794 700748 318800 700800
rect 318852 700788 318858 700800
rect 413646 700788 413652 700800
rect 318852 700760 413652 700788
rect 318852 700748 318858 700760
rect 413646 700748 413652 700760
rect 413704 700748 413710 700800
rect 218974 700680 218980 700732
rect 219032 700720 219038 700732
rect 332594 700720 332600 700732
rect 219032 700692 332600 700720
rect 219032 700680 219038 700692
rect 332594 700680 332600 700692
rect 332652 700680 332658 700732
rect 314654 700612 314660 700664
rect 314712 700652 314718 700664
rect 478506 700652 478512 700664
rect 314712 700624 478512 700652
rect 314712 700612 314718 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 154114 700544 154120 700596
rect 154172 700584 154178 700596
rect 338114 700584 338120 700596
rect 154172 700556 338120 700584
rect 154172 700544 154178 700556
rect 338114 700544 338120 700556
rect 338172 700544 338178 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 342254 700516 342260 700528
rect 89220 700488 342260 700516
rect 89220 700476 89226 700488
rect 342254 700476 342260 700488
rect 342312 700476 342318 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 340874 700448 340880 700460
rect 73028 700420 340880 700448
rect 73028 700408 73034 700420
rect 340874 700408 340880 700420
rect 340932 700408 340938 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 347866 700380 347872 700392
rect 24360 700352 347872 700380
rect 24360 700340 24366 700352
rect 347866 700340 347872 700352
rect 347924 700340 347930 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 478138 700272 478144 700324
rect 478196 700312 478202 700324
rect 559650 700312 559656 700324
rect 478196 700284 559656 700312
rect 478196 700272 478202 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 235166 698912 235172 698964
rect 235224 698952 235230 698964
rect 329834 698952 329840 698964
rect 235224 698924 329840 698952
rect 235224 698912 235230 698924
rect 329834 698912 329840 698924
rect 329892 698912 329898 698964
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 303614 696940 303620 696992
rect 303672 696980 303678 696992
rect 580166 696980 580172 696992
rect 303672 696952 580172 696980
rect 303672 696940 303678 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 304994 683136 305000 683188
rect 305052 683176 305058 683188
rect 580166 683176 580172 683188
rect 305052 683148 580172 683176
rect 305052 683136 305058 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 300854 670760 300860 670812
rect 300912 670800 300918 670812
rect 580166 670800 580172 670812
rect 300912 670772 580172 670800
rect 300912 670760 300918 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 351914 670732 351920 670744
rect 3568 670704 351920 670732
rect 3568 670692 3574 670704
rect 351914 670692 351920 670704
rect 351972 670692 351978 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 350534 656928 350540 656940
rect 3568 656900 350540 656928
rect 3568 656888 3574 656900
rect 350534 656888 350540 656900
rect 350592 656888 350598 656940
rect 298094 643084 298100 643136
rect 298152 643124 298158 643136
rect 580166 643124 580172 643136
rect 298152 643096 580172 643124
rect 298152 643084 298158 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 580166 630680 580172 630692
rect 299624 630652 580172 630680
rect 299624 630640 299630 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3326 618264 3332 618316
rect 3384 618304 3390 618316
rect 356054 618304 356060 618316
rect 3384 618276 356060 618304
rect 3384 618264 3390 618276
rect 356054 618264 356060 618276
rect 356112 618264 356118 618316
rect 296714 616836 296720 616888
rect 296772 616876 296778 616888
rect 580166 616876 580172 616888
rect 296772 616848 580172 616876
rect 296772 616836 296778 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 354674 605860 354680 605872
rect 3384 605832 354680 605860
rect 3384 605820 3390 605832
rect 354674 605820 354680 605832
rect 354732 605820 354738 605872
rect 293954 590656 293960 590708
rect 294012 590696 294018 590708
rect 579798 590696 579804 590708
rect 294012 590668 579804 590696
rect 294012 590656 294018 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 295334 576852 295340 576904
rect 295392 576892 295398 576904
rect 580166 576892 580172 576904
rect 295392 576864 580172 576892
rect 295392 576852 295398 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 361574 565876 361580 565888
rect 3108 565848 361580 565876
rect 3108 565836 3114 565848
rect 361574 565836 361580 565848
rect 361632 565836 361638 565888
rect 292574 563048 292580 563100
rect 292632 563088 292638 563100
rect 579798 563088 579804 563100
rect 292632 563060 579804 563088
rect 292632 563048 292638 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 360194 553432 360200 553444
rect 3384 553404 360200 553432
rect 3384 553392 3390 553404
rect 360194 553392 360200 553404
rect 360252 553392 360258 553444
rect 288434 536800 288440 536852
rect 288492 536840 288498 536852
rect 580166 536840 580172 536852
rect 288492 536812 580172 536840
rect 288492 536800 288498 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 289814 524424 289820 524476
rect 289872 524464 289878 524476
rect 580166 524464 580172 524476
rect 289872 524436 580172 524464
rect 289872 524424 289878 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 365714 514808 365720 514820
rect 3384 514780 365720 514808
rect 3384 514768 3390 514780
rect 365714 514768 365720 514780
rect 365772 514768 365778 514820
rect 287054 510620 287060 510672
rect 287112 510660 287118 510672
rect 580166 510660 580172 510672
rect 287112 510632 580172 510660
rect 287112 510620 287118 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 320174 502936 320180 502988
rect 320232 502976 320238 502988
rect 364334 502976 364340 502988
rect 320232 502948 364340 502976
rect 320232 502936 320238 502948
rect 364334 502936 364340 502948
rect 364392 502936 364398 502988
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 364334 501004 364340 501016
rect 3292 500976 364340 501004
rect 3292 500964 3298 500976
rect 364334 500964 364340 500976
rect 364392 500964 364398 501016
rect 284294 484372 284300 484424
rect 284352 484412 284358 484424
rect 580166 484412 580172 484424
rect 284352 484384 580172 484412
rect 284352 484372 284358 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 285858 470568 285864 470620
rect 285916 470608 285922 470620
rect 579982 470608 579988 470620
rect 285916 470580 579988 470608
rect 285916 470568 285922 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 169754 468460 169760 468512
rect 169812 468500 169818 468512
rect 334802 468500 334808 468512
rect 169812 468472 334808 468500
rect 169812 468460 169818 468472
rect 334802 468460 334808 468472
rect 334860 468460 334866 468512
rect 299474 467100 299480 467152
rect 299532 467140 299538 467152
rect 325694 467140 325700 467152
rect 299532 467112 325700 467140
rect 299532 467100 299538 467112
rect 325694 467100 325700 467112
rect 325752 467100 325758 467152
rect 316034 465672 316040 465724
rect 316092 465712 316098 465724
rect 429194 465712 429200 465724
rect 316092 465684 429200 465712
rect 316092 465672 316098 465684
rect 429194 465672 429200 465684
rect 429252 465672 429258 465724
rect 311158 464312 311164 464364
rect 311216 464352 311222 464364
rect 494054 464352 494060 464364
rect 311216 464324 494060 464352
rect 311216 464312 311222 464324
rect 494054 464312 494060 464324
rect 494112 464312 494118 464364
rect 226978 462476 226984 462528
rect 227036 462516 227042 462528
rect 375926 462516 375932 462528
rect 227036 462488 375932 462516
rect 227036 462476 227042 462488
rect 375926 462476 375932 462488
rect 375984 462476 375990 462528
rect 277118 462408 277124 462460
rect 277176 462448 277182 462460
rect 425698 462448 425704 462460
rect 277176 462420 425704 462448
rect 277176 462408 277182 462420
rect 425698 462408 425704 462420
rect 425756 462408 425762 462460
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 371234 462380 371240 462392
rect 3568 462352 371240 462380
rect 3568 462340 3574 462352
rect 371234 462340 371240 462352
rect 371292 462340 371298 462392
rect 307110 461592 307116 461644
rect 307168 461632 307174 461644
rect 478138 461632 478144 461644
rect 307168 461604 478144 461632
rect 307168 461592 307174 461604
rect 478138 461592 478144 461604
rect 478196 461592 478202 461644
rect 233970 461320 233976 461372
rect 234028 461360 234034 461372
rect 369854 461360 369860 461372
rect 234028 461332 369860 461360
rect 234028 461320 234034 461332
rect 369854 461320 369860 461332
rect 369912 461320 369918 461372
rect 280062 461252 280068 461304
rect 280120 461292 280126 461304
rect 417510 461292 417516 461304
rect 280120 461264 417516 461292
rect 280120 461252 280126 461264
rect 417510 461252 417516 461264
rect 417568 461252 417574 461304
rect 278682 461184 278688 461236
rect 278740 461224 278746 461236
rect 422938 461224 422944 461236
rect 278740 461196 422944 461224
rect 278740 461184 278746 461196
rect 422938 461184 422944 461196
rect 422996 461184 423002 461236
rect 273990 461116 273996 461168
rect 274048 461156 274054 461168
rect 421558 461156 421564 461168
rect 274048 461128 421564 461156
rect 274048 461116 274054 461128
rect 421558 461116 421564 461128
rect 421616 461116 421622 461168
rect 228358 461048 228364 461100
rect 228416 461088 228422 461100
rect 379146 461088 379152 461100
rect 228416 461060 379152 461088
rect 228416 461048 228422 461060
rect 379146 461048 379152 461060
rect 379204 461048 379210 461100
rect 229738 460980 229744 461032
rect 229796 461020 229802 461032
rect 396534 461020 396540 461032
rect 229796 460992 396540 461020
rect 229796 460980 229802 460992
rect 396534 460980 396540 460992
rect 396592 460980 396598 461032
rect 4890 460912 4896 460964
rect 4948 460952 4954 460964
rect 391934 460952 391940 460964
rect 4948 460924 391940 460952
rect 4948 460912 4954 460924
rect 391934 460912 391940 460924
rect 391992 460912 391998 460964
rect 318150 460844 318156 460896
rect 318208 460884 318214 460896
rect 397454 460884 397460 460896
rect 318208 460856 397460 460884
rect 318208 460844 318214 460856
rect 397454 460844 397460 460856
rect 397512 460844 397518 460896
rect 201494 460776 201500 460828
rect 201552 460816 201558 460828
rect 331766 460816 331772 460828
rect 201552 460788 331772 460816
rect 201552 460776 201558 460788
rect 331766 460776 331772 460788
rect 331824 460776 331830 460828
rect 313090 460708 313096 460760
rect 313148 460748 313154 460760
rect 462314 460748 462320 460760
rect 313148 460720 462320 460748
rect 313148 460708 313154 460720
rect 462314 460708 462320 460720
rect 462372 460708 462378 460760
rect 136634 460640 136640 460692
rect 136692 460680 136698 460692
rect 336734 460680 336740 460692
rect 136692 460652 336740 460680
rect 136692 460640 136698 460652
rect 336734 460640 336740 460652
rect 336792 460640 336798 460692
rect 308674 460572 308680 460624
rect 308732 460612 308738 460624
rect 527174 460612 527180 460624
rect 308732 460584 527180 460612
rect 308732 460572 308738 460584
rect 527174 460572 527180 460584
rect 527232 460572 527238 460624
rect 310238 460504 310244 460556
rect 310296 460544 310302 460556
rect 542354 460544 542360 460556
rect 310296 460516 542360 460544
rect 310296 460504 310302 460516
rect 542354 460504 542360 460516
rect 542412 460504 542418 460556
rect 104894 460436 104900 460488
rect 104952 460476 104958 460488
rect 339678 460476 339684 460488
rect 104952 460448 339684 460476
rect 104952 460436 104958 460448
rect 339678 460436 339684 460448
rect 339736 460436 339742 460488
rect 3602 460368 3608 460420
rect 3660 460408 3666 460420
rect 353846 460408 353852 460420
rect 3660 460380 353852 460408
rect 3660 460368 3666 460380
rect 353846 460368 353852 460380
rect 353904 460368 353910 460420
rect 3694 460300 3700 460352
rect 3752 460340 3758 460352
rect 358814 460340 358820 460352
rect 3752 460312 358820 460340
rect 3752 460300 3758 460312
rect 358814 460300 358820 460312
rect 358872 460300 358878 460352
rect 3786 460232 3792 460284
rect 3844 460272 3850 460284
rect 363322 460272 363328 460284
rect 3844 460244 363328 460272
rect 3844 460232 3850 460244
rect 363322 460232 363328 460244
rect 363380 460232 363386 460284
rect 3878 460164 3884 460216
rect 3936 460204 3942 460216
rect 368106 460204 368112 460216
rect 3936 460176 368112 460204
rect 3936 460164 3942 460176
rect 368106 460164 368112 460176
rect 368164 460164 368170 460216
rect 266354 460096 266360 460148
rect 266412 460136 266418 460148
rect 327074 460136 327080 460148
rect 266412 460108 327080 460136
rect 266412 460096 266418 460108
rect 327074 460096 327080 460108
rect 327132 460096 327138 460148
rect 324130 460028 324136 460080
rect 324188 460068 324194 460080
rect 347774 460068 347780 460080
rect 324188 460040 347780 460068
rect 324188 460028 324194 460040
rect 347774 460028 347780 460040
rect 347832 460028 347838 460080
rect 322842 459960 322848 460012
rect 322900 460000 322906 460012
rect 331214 460000 331220 460012
rect 322900 459972 331220 460000
rect 322900 459960 322906 459972
rect 331214 459960 331220 459972
rect 331272 459960 331278 460012
rect 349798 459620 349804 459672
rect 349856 459660 349862 459672
rect 374362 459660 374368 459672
rect 349856 459632 374368 459660
rect 349856 459620 349862 459632
rect 374362 459620 374368 459632
rect 374420 459620 374426 459672
rect 349062 459552 349068 459604
rect 349120 459592 349126 459604
rect 380894 459592 380900 459604
rect 349120 459564 380900 459592
rect 349120 459552 349126 459564
rect 380894 459552 380900 459564
rect 380952 459552 380958 459604
rect 3418 458804 3424 458856
rect 3476 458844 3482 458856
rect 349062 458844 349068 458856
rect 3476 458816 349068 458844
rect 3476 458804 3482 458816
rect 349062 458804 349068 458816
rect 349120 458804 349126 458856
rect 233878 458736 233884 458788
rect 233936 458776 233942 458788
rect 377582 458776 377588 458788
rect 233936 458748 377588 458776
rect 233936 458736 233942 458748
rect 377582 458736 377588 458748
rect 377640 458736 377646 458788
rect 275554 458668 275560 458720
rect 275612 458708 275618 458720
rect 424318 458708 424324 458720
rect 275612 458680 424324 458708
rect 275612 458668 275618 458680
rect 424318 458668 424324 458680
rect 424376 458668 424382 458720
rect 232498 458600 232504 458652
rect 232556 458640 232562 458652
rect 382274 458640 382280 458652
rect 232556 458612 382280 458640
rect 232556 458600 232562 458612
rect 382274 458600 382280 458612
rect 382332 458600 382338 458652
rect 231210 458532 231216 458584
rect 231268 458572 231274 458584
rect 387058 458572 387064 458584
rect 231268 458544 387064 458572
rect 231268 458532 231274 458544
rect 387058 458532 387064 458544
rect 387116 458532 387122 458584
rect 255038 458464 255044 458516
rect 255096 458504 255102 458516
rect 420178 458504 420184 458516
rect 255096 458476 420184 458504
rect 255096 458464 255102 458476
rect 420178 458464 420184 458476
rect 420236 458464 420242 458516
rect 245562 458396 245568 458448
rect 245620 458436 245626 458448
rect 418798 458436 418804 458448
rect 245620 458408 418804 458436
rect 245620 458396 245626 458408
rect 418798 458396 418804 458408
rect 418856 458396 418862 458448
rect 240778 458328 240784 458380
rect 240836 458368 240842 458380
rect 417418 458368 417424 458380
rect 240836 458340 417424 458368
rect 240836 458328 240842 458340
rect 417418 458328 417424 458340
rect 417476 458328 417482 458380
rect 235902 458260 235908 458312
rect 235960 458300 235966 458312
rect 580258 458300 580264 458312
rect 235960 458272 580264 458300
rect 235960 458260 235966 458272
rect 580258 458260 580264 458272
rect 580316 458260 580322 458312
rect 3602 458192 3608 458244
rect 3660 458232 3666 458244
rect 373120 458232 373126 458244
rect 3660 458204 373126 458232
rect 3660 458192 3666 458204
rect 373120 458192 373126 458204
rect 373178 458192 373184 458244
rect 273226 457660 292574 457688
rect 3510 457444 3516 457496
rect 3568 457484 3574 457496
rect 273226 457484 273254 457660
rect 281626 457580 281632 457632
rect 281684 457620 281690 457632
rect 281684 457592 287836 457620
rect 281684 457580 281690 457592
rect 3568 457456 273254 457484
rect 3568 457444 3574 457456
rect 283374 457444 283380 457496
rect 283432 457444 283438 457496
rect 283392 456804 283420 457444
rect 287808 457416 287836 457592
rect 292546 457484 292574 457660
rect 349798 457484 349804 457496
rect 292546 457456 349804 457484
rect 349798 457444 349804 457456
rect 349856 457444 349862 457496
rect 287808 457388 296714 457416
rect 296686 456872 296714 457388
rect 427078 456872 427084 456884
rect 296686 456844 427084 456872
rect 427078 456832 427084 456844
rect 427136 456832 427142 456884
rect 580166 456804 580172 456816
rect 283392 456776 580172 456804
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 233970 449868 233976 449880
rect 3384 449840 233976 449868
rect 3384 449828 3390 449840
rect 233970 449828 233976 449840
rect 234028 449828 234034 449880
rect 417510 431876 417516 431928
rect 417568 431916 417574 431928
rect 580166 431916 580172 431928
rect 417568 431888 580172 431916
rect 417568 431876 417574 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 427078 419432 427084 419484
rect 427136 419472 427142 419484
rect 580166 419472 580172 419484
rect 427136 419444 580172 419472
rect 427136 419432 427142 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 226978 411244 226984 411256
rect 3016 411216 226984 411244
rect 3016 411204 3022 411216
rect 226978 411204 226984 411216
rect 227036 411204 227042 411256
rect 422938 405628 422944 405680
rect 422996 405668 423002 405680
rect 579614 405668 579620 405680
rect 422996 405640 579620 405668
rect 422996 405628 423002 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 424318 379448 424324 379500
rect 424376 379488 424382 379500
rect 580166 379488 580172 379500
rect 424376 379460 580172 379488
rect 424376 379448 424382 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3510 372512 3516 372564
rect 3568 372552 3574 372564
rect 233878 372552 233884 372564
rect 3568 372524 233884 372552
rect 3568 372512 3574 372524
rect 233878 372512 233884 372524
rect 233936 372512 233942 372564
rect 425698 365644 425704 365696
rect 425756 365684 425762 365696
rect 580166 365684 580172 365696
rect 425756 365656 580172 365684
rect 425756 365644 425762 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 421558 353200 421564 353252
rect 421616 353240 421622 353252
rect 580166 353240 580172 353252
rect 421616 353212 580172 353240
rect 421616 353200 421622 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 228358 346372 228364 346384
rect 3200 346344 228364 346372
rect 3200 346332 3206 346344
rect 228358 346332 228364 346344
rect 228416 346332 228422 346384
rect 270540 337764 270546 337816
rect 270598 337804 270604 337816
rect 270770 337804 270776 337816
rect 270598 337776 270776 337804
rect 270598 337764 270604 337776
rect 270770 337764 270776 337776
rect 270828 337764 270834 337816
rect 331214 336880 331220 336932
rect 331272 336920 331278 336932
rect 331582 336920 331588 336932
rect 331272 336892 331588 336920
rect 331272 336880 331278 336892
rect 331582 336880 331588 336892
rect 331640 336880 331646 336932
rect 294414 336744 294420 336796
rect 294472 336744 294478 336796
rect 399018 336744 399024 336796
rect 399076 336744 399082 336796
rect 242986 336676 242992 336728
rect 243044 336716 243050 336728
rect 243262 336716 243268 336728
rect 243044 336688 243268 336716
rect 243044 336676 243050 336688
rect 243262 336676 243268 336688
rect 243320 336676 243326 336728
rect 246298 336676 246304 336728
rect 246356 336716 246362 336728
rect 247218 336716 247224 336728
rect 246356 336688 247224 336716
rect 246356 336676 246362 336688
rect 247218 336676 247224 336688
rect 247276 336676 247282 336728
rect 251818 336676 251824 336728
rect 251876 336716 251882 336728
rect 254210 336716 254216 336728
rect 251876 336688 254216 336716
rect 251876 336676 251882 336688
rect 254210 336676 254216 336688
rect 254268 336676 254274 336728
rect 269758 336676 269764 336728
rect 269816 336716 269822 336728
rect 273530 336716 273536 336728
rect 269816 336688 273536 336716
rect 269816 336676 269822 336688
rect 273530 336676 273536 336688
rect 273588 336676 273594 336728
rect 282822 336676 282828 336728
rect 282880 336716 282886 336728
rect 285674 336716 285680 336728
rect 282880 336688 285680 336716
rect 282880 336676 282886 336688
rect 285674 336676 285680 336688
rect 285732 336676 285738 336728
rect 287698 336676 287704 336728
rect 287756 336716 287762 336728
rect 290366 336716 290372 336728
rect 287756 336688 290372 336716
rect 287756 336676 287762 336688
rect 290366 336676 290372 336688
rect 290424 336676 290430 336728
rect 293218 336676 293224 336728
rect 293276 336716 293282 336728
rect 294432 336716 294460 336744
rect 293276 336688 294460 336716
rect 293276 336676 293282 336688
rect 300762 336676 300768 336728
rect 300820 336716 300826 336728
rect 304074 336716 304080 336728
rect 300820 336688 304080 336716
rect 300820 336676 300826 336688
rect 304074 336676 304080 336688
rect 304132 336676 304138 336728
rect 307018 336676 307024 336728
rect 307076 336716 307082 336728
rect 313366 336716 313372 336728
rect 307076 336688 313372 336716
rect 307076 336676 307082 336688
rect 313366 336676 313372 336688
rect 313424 336676 313430 336728
rect 316126 336676 316132 336728
rect 316184 336716 316190 336728
rect 316310 336716 316316 336728
rect 316184 336688 316316 336716
rect 316184 336676 316190 336688
rect 316310 336676 316316 336688
rect 316368 336676 316374 336728
rect 342438 336676 342444 336728
rect 342496 336716 342502 336728
rect 342622 336716 342628 336728
rect 342496 336688 342628 336716
rect 342496 336676 342502 336688
rect 342622 336676 342628 336688
rect 342680 336676 342686 336728
rect 346394 336676 346400 336728
rect 346452 336716 346458 336728
rect 346670 336716 346676 336728
rect 346452 336688 346676 336716
rect 346452 336676 346458 336688
rect 346670 336676 346676 336688
rect 346728 336676 346734 336728
rect 367094 336676 367100 336728
rect 367152 336716 367158 336728
rect 367462 336716 367468 336728
rect 367152 336688 367468 336716
rect 367152 336676 367158 336688
rect 367462 336676 367468 336688
rect 367520 336676 367526 336728
rect 386414 336676 386420 336728
rect 386472 336716 386478 336728
rect 386782 336716 386788 336728
rect 386472 336688 386788 336716
rect 386472 336676 386478 336688
rect 386782 336676 386788 336688
rect 386840 336676 386846 336728
rect 291930 336608 291936 336660
rect 291988 336648 291994 336660
rect 293310 336648 293316 336660
rect 291988 336620 293316 336648
rect 291988 336608 291994 336620
rect 293310 336608 293316 336620
rect 293368 336608 293374 336660
rect 298738 336648 298744 336660
rect 294616 336620 298744 336648
rect 294616 336592 294644 336620
rect 298738 336608 298744 336620
rect 298796 336608 298802 336660
rect 307110 336608 307116 336660
rect 307168 336648 307174 336660
rect 314838 336648 314844 336660
rect 307168 336620 314844 336648
rect 307168 336608 307174 336620
rect 314838 336608 314844 336620
rect 314896 336608 314902 336660
rect 244918 336540 244924 336592
rect 244976 336580 244982 336592
rect 246206 336580 246212 336592
rect 244976 336552 246212 336580
rect 244976 336540 244982 336552
rect 246206 336540 246212 336552
rect 246264 336540 246270 336592
rect 294598 336540 294604 336592
rect 294656 336540 294662 336592
rect 340782 336540 340788 336592
rect 340840 336580 340846 336592
rect 341334 336580 341340 336592
rect 340840 336552 341340 336580
rect 340840 336540 340846 336552
rect 341334 336540 341340 336552
rect 341392 336540 341398 336592
rect 399036 336580 399064 336744
rect 401594 336676 401600 336728
rect 401652 336716 401658 336728
rect 401870 336716 401876 336728
rect 401652 336688 401876 336716
rect 401652 336676 401658 336688
rect 401870 336676 401876 336688
rect 401928 336676 401934 336728
rect 400858 336580 400864 336592
rect 399036 336552 400864 336580
rect 400858 336540 400864 336552
rect 400916 336540 400922 336592
rect 298738 336472 298744 336524
rect 298796 336512 298802 336524
rect 302418 336512 302424 336524
rect 298796 336484 302424 336512
rect 298796 336472 298802 336484
rect 302418 336472 302424 336484
rect 302476 336472 302482 336524
rect 302970 336472 302976 336524
rect 303028 336512 303034 336524
rect 309686 336512 309692 336524
rect 303028 336484 309692 336512
rect 303028 336472 303034 336484
rect 309686 336472 309692 336484
rect 309744 336472 309750 336524
rect 350074 336472 350080 336524
rect 350132 336512 350138 336524
rect 358078 336512 358084 336524
rect 350132 336484 358084 336512
rect 350132 336472 350138 336484
rect 358078 336472 358084 336484
rect 358136 336472 358142 336524
rect 362862 336472 362868 336524
rect 362920 336512 362926 336524
rect 373350 336512 373356 336524
rect 362920 336484 373356 336512
rect 362920 336472 362926 336484
rect 373350 336472 373356 336484
rect 373408 336472 373414 336524
rect 353754 336404 353760 336456
rect 353812 336444 353818 336456
rect 382918 336444 382924 336456
rect 353812 336416 382924 336444
rect 353812 336404 353818 336416
rect 382918 336404 382924 336416
rect 382976 336404 382982 336456
rect 402330 336404 402336 336456
rect 402388 336444 402394 336456
rect 417510 336444 417516 336456
rect 402388 336416 417516 336444
rect 402388 336404 402394 336416
rect 417510 336404 417516 336416
rect 417568 336404 417574 336456
rect 231118 336336 231124 336388
rect 231176 336376 231182 336388
rect 274266 336376 274272 336388
rect 231176 336348 274272 336376
rect 231176 336336 231182 336348
rect 274266 336336 274272 336348
rect 274324 336336 274330 336388
rect 358170 336336 358176 336388
rect 358228 336376 358234 336388
rect 387058 336376 387064 336388
rect 358228 336348 387064 336376
rect 358228 336336 358234 336348
rect 387058 336336 387064 336348
rect 387116 336336 387122 336388
rect 396442 336336 396448 336388
rect 396500 336376 396506 336388
rect 424318 336376 424324 336388
rect 396500 336348 424324 336376
rect 396500 336336 396506 336348
rect 424318 336336 424324 336348
rect 424376 336336 424382 336388
rect 228358 336268 228364 336320
rect 228416 336308 228422 336320
rect 302234 336308 302240 336320
rect 228416 336280 302240 336308
rect 228416 336268 228422 336280
rect 302234 336268 302240 336280
rect 302292 336268 302298 336320
rect 315298 336268 315304 336320
rect 315356 336308 315362 336320
rect 324314 336308 324320 336320
rect 315356 336280 324320 336308
rect 315356 336268 315362 336280
rect 324314 336268 324320 336280
rect 324372 336268 324378 336320
rect 334342 336268 334348 336320
rect 334400 336308 334406 336320
rect 338206 336308 338212 336320
rect 334400 336280 338212 336308
rect 334400 336268 334406 336280
rect 338206 336268 338212 336280
rect 338264 336268 338270 336320
rect 345658 336268 345664 336320
rect 345716 336308 345722 336320
rect 357434 336308 357440 336320
rect 345716 336280 357440 336308
rect 345716 336268 345722 336280
rect 357434 336268 357440 336280
rect 357492 336268 357498 336320
rect 362770 336268 362776 336320
rect 362828 336308 362834 336320
rect 370498 336308 370504 336320
rect 362828 336280 370504 336308
rect 362828 336268 362834 336280
rect 370498 336268 370504 336280
rect 370556 336268 370562 336320
rect 373074 336268 373080 336320
rect 373132 336308 373138 336320
rect 447134 336308 447140 336320
rect 373132 336280 447140 336308
rect 373132 336268 373138 336280
rect 447134 336268 447140 336280
rect 447192 336268 447198 336320
rect 117314 336200 117320 336252
rect 117372 336240 117378 336252
rect 271046 336240 271052 336252
rect 117372 336212 271052 336240
rect 117372 336200 117378 336212
rect 271046 336200 271052 336212
rect 271104 336200 271110 336252
rect 276658 336200 276664 336252
rect 276716 336240 276722 336252
rect 277946 336240 277952 336252
rect 276716 336212 277952 336240
rect 276716 336200 276722 336212
rect 277946 336200 277952 336212
rect 278004 336200 278010 336252
rect 302878 336200 302884 336252
rect 302936 336240 302942 336252
rect 316678 336240 316684 336252
rect 302936 336212 316684 336240
rect 302936 336200 302942 336212
rect 316678 336200 316684 336212
rect 316736 336200 316742 336252
rect 339494 336200 339500 336252
rect 339552 336240 339558 336252
rect 339678 336240 339684 336252
rect 339552 336212 339684 336240
rect 339552 336200 339558 336212
rect 339678 336200 339684 336212
rect 339736 336200 339742 336252
rect 347314 336200 347320 336252
rect 347372 336240 347378 336252
rect 362954 336240 362960 336252
rect 347372 336212 362960 336240
rect 347372 336200 347378 336212
rect 362954 336200 362960 336212
rect 363012 336200 363018 336252
rect 375282 336200 375288 336252
rect 375340 336240 375346 336252
rect 454034 336240 454040 336252
rect 375340 336212 454040 336240
rect 375340 336200 375346 336212
rect 454034 336200 454040 336212
rect 454092 336200 454098 336252
rect 110414 336132 110420 336184
rect 110472 336172 110478 336184
rect 268838 336172 268844 336184
rect 110472 336144 268844 336172
rect 110472 336132 110478 336144
rect 268838 336132 268844 336144
rect 268896 336132 268902 336184
rect 297358 336132 297364 336184
rect 297416 336172 297422 336184
rect 311894 336172 311900 336184
rect 297416 336144 311900 336172
rect 297416 336132 297422 336144
rect 311894 336132 311900 336144
rect 311952 336132 311958 336184
rect 324314 336132 324320 336184
rect 324372 336172 324378 336184
rect 334894 336172 334900 336184
rect 324372 336144 334900 336172
rect 324372 336132 324378 336144
rect 334894 336132 334900 336144
rect 334952 336132 334958 336184
rect 343818 336132 343824 336184
rect 343876 336172 343882 336184
rect 345658 336172 345664 336184
rect 343876 336144 345664 336172
rect 343876 336132 343882 336144
rect 345658 336132 345664 336144
rect 345716 336132 345722 336184
rect 348602 336132 348608 336184
rect 348660 336172 348666 336184
rect 366266 336172 366272 336184
rect 348660 336144 366272 336172
rect 348660 336132 348666 336144
rect 366266 336132 366272 336144
rect 366324 336132 366330 336184
rect 377214 336132 377220 336184
rect 377272 336172 377278 336184
rect 460934 336172 460940 336184
rect 377272 336144 460940 336172
rect 377272 336132 377278 336144
rect 460934 336132 460940 336144
rect 460992 336132 460998 336184
rect 102134 336064 102140 336116
rect 102192 336104 102198 336116
rect 102192 336076 258074 336104
rect 102192 336064 102198 336076
rect 10318 335996 10324 336048
rect 10376 336036 10382 336048
rect 236638 336036 236644 336048
rect 10376 336008 236644 336036
rect 10376 335996 10382 336008
rect 236638 335996 236644 336008
rect 236696 335996 236702 336048
rect 258046 336036 258074 336076
rect 264238 336064 264244 336116
rect 264296 336104 264302 336116
rect 264974 336104 264980 336116
rect 264296 336076 264980 336104
rect 264296 336064 264302 336076
rect 264974 336064 264980 336076
rect 265032 336064 265038 336116
rect 289078 336064 289084 336116
rect 289136 336104 289142 336116
rect 310790 336104 310796 336116
rect 289136 336076 310796 336104
rect 289136 336064 289142 336076
rect 310790 336064 310796 336076
rect 310848 336064 310854 336116
rect 318058 336064 318064 336116
rect 318116 336104 318122 336116
rect 331214 336104 331220 336116
rect 318116 336076 331220 336104
rect 318116 336064 318122 336076
rect 331214 336064 331220 336076
rect 331272 336064 331278 336116
rect 350810 336064 350816 336116
rect 350868 336104 350874 336116
rect 373994 336104 374000 336116
rect 350868 336076 374000 336104
rect 350868 336064 350874 336076
rect 373994 336064 374000 336076
rect 374052 336064 374058 336116
rect 379882 336064 379888 336116
rect 379940 336104 379946 336116
rect 467834 336104 467840 336116
rect 379940 336076 467840 336104
rect 379940 336064 379946 336076
rect 467834 336064 467840 336076
rect 467892 336064 467898 336116
rect 266722 336036 266728 336048
rect 258046 336008 266728 336036
rect 266722 335996 266728 336008
rect 266780 335996 266786 336048
rect 276750 335996 276756 336048
rect 276808 336036 276814 336048
rect 284478 336036 284484 336048
rect 276808 336008 284484 336036
rect 276808 335996 276814 336008
rect 284478 335996 284484 336008
rect 284536 335996 284542 336048
rect 286226 335996 286232 336048
rect 286284 336036 286290 336048
rect 291194 336036 291200 336048
rect 286284 336008 291200 336036
rect 286284 335996 286290 336008
rect 291194 335996 291200 336008
rect 291252 335996 291258 336048
rect 291838 335996 291844 336048
rect 291896 336036 291902 336048
rect 315206 336036 315212 336048
rect 291896 336008 315212 336036
rect 291896 335996 291902 336008
rect 315206 335996 315212 336008
rect 315264 335996 315270 336048
rect 320174 335996 320180 336048
rect 320232 336036 320238 336048
rect 333974 336036 333980 336048
rect 320232 336008 333980 336036
rect 320232 335996 320238 336008
rect 333974 335996 333980 336008
rect 334032 335996 334038 336048
rect 344922 335996 344928 336048
rect 344980 336036 344986 336048
rect 351178 336036 351184 336048
rect 344980 336008 351184 336036
rect 344980 335996 344986 336008
rect 351178 335996 351184 336008
rect 351236 335996 351242 336048
rect 351914 335996 351920 336048
rect 351972 336036 351978 336048
rect 377398 336036 377404 336048
rect 351972 336008 377404 336036
rect 351972 335996 351978 336008
rect 377398 335996 377404 336008
rect 377456 335996 377462 336048
rect 381814 335996 381820 336048
rect 381872 336036 381878 336048
rect 474734 336036 474740 336048
rect 381872 336008 474740 336036
rect 381872 335996 381878 336008
rect 474734 335996 474740 336008
rect 474792 335996 474798 336048
rect 260834 335928 260840 335980
rect 260892 335968 260898 335980
rect 261110 335968 261116 335980
rect 260892 335940 261116 335968
rect 260892 335928 260898 335940
rect 261110 335928 261116 335940
rect 261168 335928 261174 335980
rect 305638 335928 305644 335980
rect 305696 335968 305702 335980
rect 307202 335968 307208 335980
rect 305696 335940 307208 335968
rect 305696 335928 305702 335940
rect 307202 335928 307208 335940
rect 307260 335928 307266 335980
rect 271138 335792 271144 335844
rect 271196 335832 271202 335844
rect 272426 335832 272432 335844
rect 271196 335804 272432 335832
rect 271196 335792 271202 335804
rect 272426 335792 272432 335804
rect 272484 335792 272490 335844
rect 319438 335792 319444 335844
rect 319496 335832 319502 335844
rect 321002 335832 321008 335844
rect 319496 335804 321008 335832
rect 319496 335792 319502 335804
rect 321002 335792 321008 335804
rect 321060 335792 321066 335844
rect 286410 335724 286416 335776
rect 286468 335764 286474 335776
rect 287790 335764 287796 335776
rect 286468 335736 287796 335764
rect 286468 335724 286474 335736
rect 287790 335724 287796 335736
rect 287848 335724 287854 335776
rect 320818 335724 320824 335776
rect 320876 335764 320882 335776
rect 326522 335764 326528 335776
rect 320876 335736 326528 335764
rect 320876 335724 320882 335736
rect 326522 335724 326528 335736
rect 326580 335724 326586 335776
rect 297450 335656 297456 335708
rect 297508 335696 297514 335708
rect 299842 335696 299848 335708
rect 297508 335668 299848 335696
rect 297508 335656 297514 335668
rect 299842 335656 299848 335668
rect 299900 335656 299906 335708
rect 340966 335656 340972 335708
rect 341024 335696 341030 335708
rect 342254 335696 342260 335708
rect 341024 335668 342260 335696
rect 341024 335656 341030 335668
rect 342254 335656 342260 335668
rect 342312 335656 342318 335708
rect 303522 335588 303528 335640
rect 303580 335628 303586 335640
rect 306466 335628 306472 335640
rect 303580 335600 306472 335628
rect 303580 335588 303586 335600
rect 306466 335588 306472 335600
rect 306524 335588 306530 335640
rect 289170 335520 289176 335572
rect 289228 335560 289234 335572
rect 289998 335560 290004 335572
rect 289228 335532 290004 335560
rect 289228 335520 289234 335532
rect 289998 335520 290004 335532
rect 290056 335520 290062 335572
rect 411806 335452 411812 335504
rect 411864 335492 411870 335504
rect 413278 335492 413284 335504
rect 411864 335464 413284 335492
rect 411864 335452 411870 335464
rect 413278 335452 413284 335464
rect 413336 335452 413342 335504
rect 301498 335384 301504 335436
rect 301556 335424 301562 335436
rect 308582 335424 308588 335436
rect 301556 335396 308588 335424
rect 301556 335384 301562 335396
rect 308582 335384 308588 335396
rect 308640 335384 308646 335436
rect 379974 335384 379980 335436
rect 380032 335424 380038 335436
rect 381538 335424 381544 335436
rect 380032 335396 381544 335424
rect 380032 335384 380038 335396
rect 381538 335384 381544 335396
rect 381596 335384 381602 335436
rect 233970 335316 233976 335368
rect 234028 335356 234034 335368
rect 240134 335356 240140 335368
rect 234028 335328 240140 335356
rect 234028 335316 234034 335328
rect 240134 335316 240140 335328
rect 240192 335316 240198 335368
rect 295978 335316 295984 335368
rect 296036 335356 296042 335368
rect 296714 335356 296720 335368
rect 296036 335328 296720 335356
rect 296036 335316 296042 335328
rect 296714 335316 296720 335328
rect 296772 335316 296778 335368
rect 304258 335316 304264 335368
rect 304316 335356 304322 335368
rect 307846 335356 307852 335368
rect 304316 335328 307852 335356
rect 304316 335316 304322 335328
rect 307846 335316 307852 335328
rect 307904 335316 307910 335368
rect 313918 335316 313924 335368
rect 313976 335356 313982 335368
rect 317414 335356 317420 335368
rect 313976 335328 317420 335356
rect 313976 335316 313982 335328
rect 317414 335316 317420 335328
rect 317472 335316 317478 335368
rect 331582 335316 331588 335368
rect 331640 335356 331646 335368
rect 337102 335356 337108 335368
rect 331640 335328 337108 335356
rect 331640 335316 331646 335328
rect 337102 335316 337108 335328
rect 337160 335316 337166 335368
rect 224954 334636 224960 334688
rect 225012 334676 225018 334688
rect 300762 334676 300768 334688
rect 225012 334648 300768 334676
rect 225012 334636 225018 334648
rect 300762 334636 300768 334648
rect 300820 334636 300826 334688
rect 383562 334636 383568 334688
rect 383620 334676 383626 334688
rect 480254 334676 480260 334688
rect 383620 334648 480260 334676
rect 383620 334636 383626 334648
rect 480254 334636 480260 334648
rect 480312 334636 480318 334688
rect 3418 334568 3424 334620
rect 3476 334608 3482 334620
rect 234798 334608 234804 334620
rect 3476 334580 234804 334608
rect 3476 334568 3482 334580
rect 234798 334568 234804 334580
rect 234856 334568 234862 334620
rect 405274 334568 405280 334620
rect 405332 334608 405338 334620
rect 550634 334608 550640 334620
rect 405332 334580 550640 334608
rect 405332 334568 405338 334580
rect 550634 334568 550640 334580
rect 550692 334568 550698 334620
rect 384482 333276 384488 333328
rect 384540 333316 384546 333328
rect 483014 333316 483020 333328
rect 384540 333288 483020 333316
rect 384540 333276 384546 333288
rect 483014 333276 483020 333288
rect 483072 333276 483078 333328
rect 303522 333248 303528 333260
rect 238726 333220 303528 333248
rect 231854 333140 231860 333192
rect 231912 333180 231918 333192
rect 238726 333180 238754 333220
rect 303522 333208 303528 333220
rect 303580 333208 303586 333260
rect 561674 333248 561680 333260
rect 412606 333220 561680 333248
rect 231912 333152 238754 333180
rect 231912 333140 231918 333152
rect 408586 333140 408592 333192
rect 408644 333180 408650 333192
rect 412606 333180 412634 333220
rect 561674 333208 561680 333220
rect 561732 333208 561738 333260
rect 408644 333152 412634 333180
rect 408644 333140 408650 333152
rect 175274 331916 175280 331968
rect 175332 331956 175338 331968
rect 288894 331956 288900 331968
rect 175332 331928 288900 331956
rect 175332 331916 175338 331928
rect 288894 331916 288900 331928
rect 288952 331916 288958 331968
rect 46934 331848 46940 331900
rect 46992 331888 46998 331900
rect 249426 331888 249432 331900
rect 46992 331860 249432 331888
rect 46992 331848 46998 331860
rect 249426 331848 249432 331860
rect 249484 331848 249490 331900
rect 397546 331848 397552 331900
rect 397604 331888 397610 331900
rect 525794 331888 525800 331900
rect 397604 331860 525800 331888
rect 397604 331848 397610 331860
rect 525794 331848 525800 331860
rect 525852 331848 525858 331900
rect 280430 331168 280436 331220
rect 280488 331208 280494 331220
rect 280614 331208 280620 331220
rect 280488 331180 280620 331208
rect 280488 331168 280494 331180
rect 280614 331168 280620 331180
rect 280672 331168 280678 331220
rect 283190 330760 283196 330812
rect 283248 330800 283254 330812
rect 283466 330800 283472 330812
rect 283248 330772 283472 330800
rect 283248 330760 283254 330772
rect 283466 330760 283472 330772
rect 283524 330760 283530 330812
rect 234586 330704 258074 330732
rect 168374 330556 168380 330608
rect 168432 330596 168438 330608
rect 234586 330596 234614 330704
rect 252738 330664 252744 330676
rect 168432 330568 234614 330596
rect 249628 330636 252744 330664
rect 168432 330556 168438 330568
rect 57974 330488 57980 330540
rect 58032 330528 58038 330540
rect 249628 330528 249656 330636
rect 252738 330624 252744 330636
rect 252796 330624 252802 330676
rect 258046 330596 258074 330704
rect 286686 330596 286692 330608
rect 258046 330568 286692 330596
rect 286686 330556 286692 330568
rect 286744 330556 286750 330608
rect 390002 330556 390008 330608
rect 390060 330596 390066 330608
rect 500954 330596 500960 330608
rect 390060 330568 500960 330596
rect 390060 330556 390066 330568
rect 500954 330556 500960 330568
rect 501012 330556 501018 330608
rect 58032 330500 249656 330528
rect 58032 330488 58038 330500
rect 249794 330488 249800 330540
rect 249852 330528 249858 330540
rect 250162 330528 250168 330540
rect 249852 330500 250168 330528
rect 249852 330488 249858 330500
rect 250162 330488 250168 330500
rect 250220 330488 250226 330540
rect 251174 330488 251180 330540
rect 251232 330528 251238 330540
rect 252002 330528 252008 330540
rect 251232 330500 252008 330528
rect 251232 330488 251238 330500
rect 252002 330488 252008 330500
rect 252060 330488 252066 330540
rect 254026 330488 254032 330540
rect 254084 330528 254090 330540
rect 254946 330528 254952 330540
rect 254084 330500 254952 330528
rect 254084 330488 254090 330500
rect 254946 330488 254952 330500
rect 255004 330488 255010 330540
rect 255406 330488 255412 330540
rect 255464 330528 255470 330540
rect 255682 330528 255688 330540
rect 255464 330500 255688 330528
rect 255464 330488 255470 330500
rect 255682 330488 255688 330500
rect 255740 330488 255746 330540
rect 256694 330488 256700 330540
rect 256752 330528 256758 330540
rect 257154 330528 257160 330540
rect 256752 330500 257160 330528
rect 256752 330488 256758 330500
rect 257154 330488 257160 330500
rect 257212 330488 257218 330540
rect 258166 330488 258172 330540
rect 258224 330528 258230 330540
rect 258626 330528 258632 330540
rect 258224 330500 258632 330528
rect 258224 330488 258230 330500
rect 258626 330488 258632 330500
rect 258684 330488 258690 330540
rect 260926 330488 260932 330540
rect 260984 330528 260990 330540
rect 261846 330528 261852 330540
rect 260984 330500 261852 330528
rect 260984 330488 260990 330500
rect 261846 330488 261852 330500
rect 261904 330488 261910 330540
rect 262306 330488 262312 330540
rect 262364 330528 262370 330540
rect 263318 330528 263324 330540
rect 262364 330500 263324 330528
rect 262364 330488 262370 330500
rect 263318 330488 263324 330500
rect 263376 330488 263382 330540
rect 266538 330488 266544 330540
rect 266596 330528 266602 330540
rect 266998 330528 267004 330540
rect 266596 330500 267004 330528
rect 266596 330488 266602 330500
rect 266998 330488 267004 330500
rect 267056 330488 267062 330540
rect 267826 330488 267832 330540
rect 267884 330528 267890 330540
rect 268470 330528 268476 330540
rect 267884 330500 268476 330528
rect 267884 330488 267890 330500
rect 268470 330488 268476 330500
rect 268528 330488 268534 330540
rect 269114 330488 269120 330540
rect 269172 330528 269178 330540
rect 269942 330528 269948 330540
rect 269172 330500 269948 330528
rect 269172 330488 269178 330500
rect 269942 330488 269948 330500
rect 270000 330488 270006 330540
rect 270586 330488 270592 330540
rect 270644 330528 270650 330540
rect 271322 330528 271328 330540
rect 270644 330500 271328 330528
rect 270644 330488 270650 330500
rect 271322 330488 271328 330500
rect 271380 330488 271386 330540
rect 271966 330488 271972 330540
rect 272024 330528 272030 330540
rect 272794 330528 272800 330540
rect 272024 330500 272800 330528
rect 272024 330488 272030 330500
rect 272794 330488 272800 330500
rect 272852 330488 272858 330540
rect 285766 330488 285772 330540
rect 285824 330528 285830 330540
rect 286318 330528 286324 330540
rect 285824 330500 286324 330528
rect 285824 330488 285830 330500
rect 286318 330488 286324 330500
rect 286376 330488 286382 330540
rect 287146 330488 287152 330540
rect 287204 330528 287210 330540
rect 288158 330528 288164 330540
rect 287204 330500 288164 330528
rect 287204 330488 287210 330500
rect 288158 330488 288164 330500
rect 288216 330488 288222 330540
rect 291378 330488 291384 330540
rect 291436 330528 291442 330540
rect 292206 330528 292212 330540
rect 291436 330500 292212 330528
rect 291436 330488 291442 330500
rect 292206 330488 292212 330500
rect 292264 330488 292270 330540
rect 294230 330488 294236 330540
rect 294288 330528 294294 330540
rect 295150 330528 295156 330540
rect 294288 330500 295156 330528
rect 294288 330488 294294 330500
rect 295150 330488 295156 330500
rect 295208 330488 295214 330540
rect 295334 330488 295340 330540
rect 295392 330528 295398 330540
rect 295794 330528 295800 330540
rect 295392 330500 295800 330528
rect 295392 330488 295398 330500
rect 295794 330488 295800 330500
rect 295852 330488 295858 330540
rect 298370 330488 298376 330540
rect 298428 330528 298434 330540
rect 299106 330528 299112 330540
rect 298428 330500 299112 330528
rect 298428 330488 298434 330500
rect 299106 330488 299112 330500
rect 299164 330488 299170 330540
rect 299566 330488 299572 330540
rect 299624 330528 299630 330540
rect 300578 330528 300584 330540
rect 299624 330500 300584 330528
rect 299624 330488 299630 330500
rect 300578 330488 300584 330500
rect 300636 330488 300642 330540
rect 300854 330488 300860 330540
rect 300912 330528 300918 330540
rect 301682 330528 301688 330540
rect 300912 330500 301688 330528
rect 300912 330488 300918 330500
rect 301682 330488 301688 330500
rect 301740 330488 301746 330540
rect 313458 330488 313464 330540
rect 313516 330528 313522 330540
rect 314102 330528 314108 330540
rect 313516 330500 314108 330528
rect 313516 330488 313522 330500
rect 314102 330488 314108 330500
rect 314160 330488 314166 330540
rect 317690 330488 317696 330540
rect 317748 330528 317754 330540
rect 318150 330528 318156 330540
rect 317748 330500 318156 330528
rect 317748 330488 317754 330500
rect 318150 330488 318156 330500
rect 318208 330488 318214 330540
rect 318794 330488 318800 330540
rect 318852 330528 318858 330540
rect 319254 330528 319260 330540
rect 318852 330500 319260 330528
rect 318852 330488 318858 330500
rect 319254 330488 319260 330500
rect 319312 330488 319318 330540
rect 332594 330488 332600 330540
rect 332652 330528 332658 330540
rect 333054 330528 333060 330540
rect 332652 330500 333060 330528
rect 332652 330488 332658 330500
rect 333054 330488 333060 330500
rect 333112 330488 333118 330540
rect 335354 330488 335360 330540
rect 335412 330528 335418 330540
rect 335998 330528 336004 330540
rect 335412 330500 336004 330528
rect 335412 330488 335418 330500
rect 335998 330488 336004 330500
rect 336056 330488 336062 330540
rect 360194 330488 360200 330540
rect 360252 330528 360258 330540
rect 360838 330528 360844 330540
rect 360252 330500 360844 330528
rect 360252 330488 360258 330500
rect 360838 330488 360844 330500
rect 360896 330488 360902 330540
rect 363138 330488 363144 330540
rect 363196 330528 363202 330540
rect 363782 330528 363788 330540
rect 363196 330500 363788 330528
rect 363196 330488 363202 330500
rect 363782 330488 363788 330500
rect 363840 330488 363846 330540
rect 364426 330488 364432 330540
rect 364484 330528 364490 330540
rect 365254 330528 365260 330540
rect 364484 330500 365260 330528
rect 364484 330488 364490 330500
rect 365254 330488 365260 330500
rect 365312 330488 365318 330540
rect 365806 330488 365812 330540
rect 365864 330528 365870 330540
rect 366726 330528 366732 330540
rect 365864 330500 366732 330528
rect 365864 330488 365870 330500
rect 366726 330488 366732 330500
rect 366784 330488 366790 330540
rect 368474 330488 368480 330540
rect 368532 330528 368538 330540
rect 369578 330528 369584 330540
rect 368532 330500 369584 330528
rect 368532 330488 368538 330500
rect 369578 330488 369584 330500
rect 369636 330488 369642 330540
rect 390738 330488 390744 330540
rect 390796 330528 390802 330540
rect 391198 330528 391204 330540
rect 390796 330500 391204 330528
rect 390796 330488 390802 330500
rect 391198 330488 391204 330500
rect 391256 330488 391262 330540
rect 392026 330488 392032 330540
rect 392084 330528 392090 330540
rect 392578 330528 392584 330540
rect 392084 330500 392584 330528
rect 392084 330488 392090 330500
rect 392578 330488 392584 330500
rect 392636 330488 392642 330540
rect 393406 330488 393412 330540
rect 393464 330528 393470 330540
rect 394418 330528 394424 330540
rect 393464 330500 394424 330528
rect 393464 330488 393470 330500
rect 394418 330488 394424 330500
rect 394476 330488 394482 330540
rect 394694 330488 394700 330540
rect 394752 330528 394758 330540
rect 395154 330528 395160 330540
rect 394752 330500 395160 330528
rect 394752 330488 394758 330500
rect 395154 330488 395160 330500
rect 395212 330488 395218 330540
rect 397454 330488 397460 330540
rect 397512 330528 397518 330540
rect 398098 330528 398104 330540
rect 397512 330500 398104 330528
rect 397512 330488 397518 330500
rect 398098 330488 398104 330500
rect 398156 330488 398162 330540
rect 408494 330488 408500 330540
rect 408552 330528 408558 330540
rect 409046 330528 409052 330540
rect 408552 330500 409052 330528
rect 408552 330488 408558 330500
rect 409046 330488 409052 330500
rect 409104 330488 409110 330540
rect 409966 330488 409972 330540
rect 410024 330528 410030 330540
rect 410886 330528 410892 330540
rect 410024 330500 410892 330528
rect 410024 330488 410030 330500
rect 410886 330488 410892 330500
rect 410944 330488 410950 330540
rect 411346 330488 411352 330540
rect 411404 330528 411410 330540
rect 412358 330528 412364 330540
rect 411404 330500 412364 330528
rect 411404 330488 411410 330500
rect 412358 330488 412364 330500
rect 412416 330488 412422 330540
rect 567194 330528 567200 330540
rect 412606 330500 567200 330528
rect 244274 330420 244280 330472
rect 244332 330460 244338 330472
rect 244734 330460 244740 330472
rect 244332 330432 244740 330460
rect 244332 330420 244338 330432
rect 244734 330420 244740 330432
rect 244792 330420 244798 330472
rect 249886 330420 249892 330472
rect 249944 330460 249950 330472
rect 250898 330460 250904 330472
rect 249944 330432 250904 330460
rect 249944 330420 249950 330432
rect 250898 330420 250904 330432
rect 250956 330420 250962 330472
rect 255314 330420 255320 330472
rect 255372 330460 255378 330472
rect 256418 330460 256424 330472
rect 255372 330432 256424 330460
rect 255372 330420 255378 330432
rect 256418 330420 256424 330432
rect 256476 330420 256482 330472
rect 256786 330420 256792 330472
rect 256844 330460 256850 330472
rect 257522 330460 257528 330472
rect 256844 330432 257528 330460
rect 256844 330420 256850 330432
rect 257522 330420 257528 330432
rect 257580 330420 257586 330472
rect 258258 330420 258264 330472
rect 258316 330460 258322 330472
rect 258994 330460 259000 330472
rect 258316 330432 259000 330460
rect 258316 330420 258322 330432
rect 258994 330420 259000 330432
rect 259052 330420 259058 330472
rect 266446 330420 266452 330472
rect 266504 330460 266510 330472
rect 267366 330460 267372 330472
rect 266504 330432 267372 330460
rect 266504 330420 266510 330432
rect 267366 330420 267372 330432
rect 267424 330420 267430 330472
rect 317506 330420 317512 330472
rect 317564 330460 317570 330472
rect 318518 330460 318524 330472
rect 317564 330432 318524 330460
rect 317564 330420 317570 330432
rect 318518 330420 318524 330432
rect 318576 330420 318582 330472
rect 318978 330420 318984 330472
rect 319036 330460 319042 330472
rect 319898 330460 319904 330472
rect 319036 330432 319904 330460
rect 319036 330420 319042 330432
rect 319898 330420 319904 330432
rect 319956 330420 319962 330472
rect 332686 330420 332692 330472
rect 332744 330460 332750 330472
rect 333422 330460 333428 330472
rect 332744 330432 333428 330460
rect 332744 330420 332750 330432
rect 333422 330420 333428 330432
rect 333480 330420 333486 330472
rect 390554 330420 390560 330472
rect 390612 330460 390618 330472
rect 391474 330460 391480 330472
rect 390612 330432 391480 330460
rect 390612 330420 390618 330432
rect 391474 330420 391480 330432
rect 391532 330420 391538 330472
rect 391934 330420 391940 330472
rect 391992 330460 391998 330472
rect 392946 330460 392952 330472
rect 391992 330432 392952 330460
rect 391992 330420 391998 330432
rect 392946 330420 392952 330432
rect 393004 330420 393010 330472
rect 410426 330420 410432 330472
rect 410484 330460 410490 330472
rect 412606 330460 412634 330500
rect 567194 330488 567200 330500
rect 567252 330488 567258 330540
rect 410484 330432 412634 330460
rect 410484 330420 410490 330432
rect 258074 330352 258080 330404
rect 258132 330392 258138 330404
rect 258442 330392 258448 330404
rect 258132 330364 258448 330392
rect 258132 330352 258138 330364
rect 258442 330352 258448 330364
rect 258500 330352 258506 330404
rect 296990 330352 296996 330404
rect 297048 330392 297054 330404
rect 297634 330392 297640 330404
rect 297048 330364 297640 330392
rect 297048 330352 297054 330364
rect 297634 330352 297640 330364
rect 297692 330352 297698 330404
rect 361574 329672 361580 329724
rect 361632 329712 361638 329724
rect 361942 329712 361948 329724
rect 361632 329684 361948 329712
rect 361632 329672 361638 329684
rect 361942 329672 361948 329684
rect 362000 329672 362006 329724
rect 396166 329672 396172 329724
rect 396224 329712 396230 329724
rect 396994 329712 397000 329724
rect 396224 329684 397000 329712
rect 396224 329672 396230 329684
rect 396994 329672 397000 329684
rect 397052 329672 397058 329724
rect 262214 329264 262220 329316
rect 262272 329304 262278 329316
rect 262950 329304 262956 329316
rect 262272 329276 262956 329304
rect 262272 329264 262278 329276
rect 262950 329264 262956 329276
rect 263008 329264 263014 329316
rect 164234 329128 164240 329180
rect 164292 329168 164298 329180
rect 282822 329168 282828 329180
rect 164292 329140 282828 329168
rect 164292 329128 164298 329140
rect 282822 329128 282828 329140
rect 282880 329128 282886 329180
rect 283006 329128 283012 329180
rect 283064 329168 283070 329180
rect 283742 329168 283748 329180
rect 283064 329140 283748 329168
rect 283064 329128 283070 329140
rect 283742 329128 283748 329140
rect 283800 329128 283806 329180
rect 60734 329060 60740 329112
rect 60792 329100 60798 329112
rect 253934 329100 253940 329112
rect 60792 329072 253940 329100
rect 60792 329060 60798 329072
rect 253934 329060 253940 329072
rect 253992 329060 253998 329112
rect 367278 329060 367284 329112
rect 367336 329100 367342 329112
rect 368106 329100 368112 329112
rect 367336 329072 368112 329100
rect 367336 329060 367342 329072
rect 368106 329060 368112 329072
rect 368164 329060 368170 329112
rect 392118 329060 392124 329112
rect 392176 329100 392182 329112
rect 507854 329100 507860 329112
rect 392176 329072 507860 329100
rect 392176 329060 392182 329072
rect 507854 329060 507860 329072
rect 507912 329060 507918 329112
rect 314838 328788 314844 328840
rect 314896 328828 314902 328840
rect 315574 328828 315580 328840
rect 314896 328800 315580 328828
rect 314896 328788 314902 328800
rect 315574 328788 315580 328800
rect 315632 328788 315638 328840
rect 295426 328720 295432 328772
rect 295484 328760 295490 328772
rect 296162 328760 296168 328772
rect 295484 328732 296168 328760
rect 295484 328720 295490 328732
rect 296162 328720 296168 328732
rect 296220 328720 296226 328772
rect 245746 328516 245752 328568
rect 245804 328556 245810 328568
rect 246574 328556 246580 328568
rect 245804 328528 246580 328556
rect 245804 328516 245810 328528
rect 246574 328516 246580 328528
rect 246632 328516 246638 328568
rect 265158 327972 265164 328024
rect 265216 328012 265222 328024
rect 265894 328012 265900 328024
rect 265216 327984 265900 328012
rect 265216 327972 265222 327984
rect 265894 327972 265900 327984
rect 265952 327972 265958 328024
rect 365714 327836 365720 327888
rect 365772 327876 365778 327888
rect 366358 327876 366364 327888
rect 365772 327848 366364 327876
rect 365772 327836 365778 327848
rect 366358 327836 366364 327848
rect 366416 327836 366422 327888
rect 201494 327768 201500 327820
rect 201552 327808 201558 327820
rect 296714 327808 296720 327820
rect 201552 327780 296720 327808
rect 201552 327768 201558 327780
rect 296714 327768 296720 327780
rect 296772 327768 296778 327820
rect 396074 327768 396080 327820
rect 396132 327808 396138 327820
rect 396626 327808 396632 327820
rect 396132 327780 396632 327808
rect 396132 327768 396138 327780
rect 396626 327768 396632 327780
rect 396684 327768 396690 327820
rect 125594 327700 125600 327752
rect 125652 327740 125658 327752
rect 269758 327740 269764 327752
rect 125652 327712 269764 327740
rect 125652 327700 125658 327712
rect 269758 327700 269764 327712
rect 269816 327700 269822 327752
rect 394050 327700 394056 327752
rect 394108 327740 394114 327752
rect 514754 327740 514760 327752
rect 394108 327712 514760 327740
rect 394108 327700 394114 327712
rect 514754 327700 514760 327712
rect 514812 327700 514818 327752
rect 259546 327632 259552 327684
rect 259604 327672 259610 327684
rect 260374 327672 260380 327684
rect 259604 327644 260380 327672
rect 259604 327632 259610 327644
rect 260374 327632 260380 327644
rect 260432 327632 260438 327684
rect 367186 327632 367192 327684
rect 367244 327672 367250 327684
rect 367738 327672 367744 327684
rect 367244 327644 367744 327672
rect 367244 327632 367250 327644
rect 367738 327632 367744 327644
rect 367796 327632 367802 327684
rect 393314 327632 393320 327684
rect 393372 327672 393378 327684
rect 393682 327672 393688 327684
rect 393372 327644 393688 327672
rect 393372 327632 393378 327644
rect 393682 327632 393688 327644
rect 393740 327632 393746 327684
rect 378318 326680 378324 326732
rect 378376 326680 378382 326732
rect 383746 326680 383752 326732
rect 383804 326720 383810 326732
rect 383804 326692 383884 326720
rect 383804 326680 383810 326692
rect 378336 326528 378364 326680
rect 383856 326528 383884 326692
rect 237558 326476 237564 326528
rect 237616 326516 237622 326528
rect 237742 326516 237748 326528
rect 237616 326488 237748 326516
rect 237616 326476 237622 326488
rect 237742 326476 237748 326488
rect 237800 326476 237806 326528
rect 241790 326476 241796 326528
rect 241848 326516 241854 326528
rect 241974 326516 241980 326528
rect 241848 326488 241980 326516
rect 241848 326476 241854 326488
rect 241974 326476 241980 326488
rect 242032 326476 242038 326528
rect 354950 326476 354956 326528
rect 355008 326516 355014 326528
rect 355134 326516 355140 326528
rect 355008 326488 355140 326516
rect 355008 326476 355014 326488
rect 355134 326476 355140 326488
rect 355192 326476 355198 326528
rect 375558 326476 375564 326528
rect 375616 326516 375622 326528
rect 375742 326516 375748 326528
rect 375616 326488 375748 326516
rect 375616 326476 375622 326488
rect 375742 326476 375748 326488
rect 375800 326476 375806 326528
rect 378318 326476 378324 326528
rect 378376 326476 378382 326528
rect 381078 326476 381084 326528
rect 381136 326516 381142 326528
rect 381262 326516 381268 326528
rect 381136 326488 381268 326516
rect 381136 326476 381142 326488
rect 381262 326476 381268 326488
rect 381320 326476 381326 326528
rect 383838 326476 383844 326528
rect 383896 326476 383902 326528
rect 193214 326408 193220 326460
rect 193272 326448 193278 326460
rect 293218 326448 293224 326460
rect 193272 326420 293224 326448
rect 193272 326408 193278 326420
rect 293218 326408 293224 326420
rect 293276 326408 293282 326460
rect 323026 326408 323032 326460
rect 323084 326448 323090 326460
rect 323946 326448 323952 326460
rect 323084 326420 323952 326448
rect 323084 326408 323090 326420
rect 323946 326408 323952 326420
rect 324004 326408 324010 326460
rect 328454 326408 328460 326460
rect 328512 326448 328518 326460
rect 329098 326448 329104 326460
rect 328512 326420 329104 326448
rect 328512 326408 328518 326420
rect 329098 326408 329104 326420
rect 329156 326408 329162 326460
rect 329926 326408 329932 326460
rect 329984 326448 329990 326460
rect 330570 326448 330576 326460
rect 329984 326420 330576 326448
rect 329984 326408 329990 326420
rect 330570 326408 330576 326420
rect 330628 326408 330634 326460
rect 354674 326408 354680 326460
rect 354732 326448 354738 326460
rect 355686 326448 355692 326460
rect 354732 326420 355692 326448
rect 354732 326408 354738 326420
rect 355686 326408 355692 326420
rect 355744 326408 355750 326460
rect 356238 326408 356244 326460
rect 356296 326448 356302 326460
rect 356422 326448 356428 326460
rect 356296 326420 356428 326448
rect 356296 326408 356302 326420
rect 356422 326408 356428 326420
rect 356480 326408 356486 326460
rect 369854 326408 369860 326460
rect 369912 326448 369918 326460
rect 370682 326448 370688 326460
rect 369912 326420 370688 326448
rect 369912 326408 369918 326420
rect 370682 326408 370688 326420
rect 370740 326408 370746 326460
rect 371418 326408 371424 326460
rect 371476 326448 371482 326460
rect 372154 326448 372160 326460
rect 371476 326420 372160 326448
rect 371476 326408 371482 326420
rect 372154 326408 372160 326420
rect 372212 326408 372218 326460
rect 372706 326408 372712 326460
rect 372764 326448 372770 326460
rect 373626 326448 373632 326460
rect 372764 326420 373632 326448
rect 372764 326408 372770 326420
rect 373626 326408 373632 326420
rect 373684 326408 373690 326460
rect 374178 326408 374184 326460
rect 374236 326448 374242 326460
rect 374730 326448 374736 326460
rect 374236 326420 374736 326448
rect 374236 326408 374242 326420
rect 374730 326408 374736 326420
rect 374788 326408 374794 326460
rect 375374 326408 375380 326460
rect 375432 326448 375438 326460
rect 376202 326448 376208 326460
rect 375432 326420 376208 326448
rect 375432 326408 375438 326420
rect 376202 326408 376208 326420
rect 376260 326408 376266 326460
rect 376846 326408 376852 326460
rect 376904 326448 376910 326460
rect 377030 326448 377036 326460
rect 376904 326420 377036 326448
rect 376904 326408 376910 326420
rect 377030 326408 377036 326420
rect 377088 326408 377094 326460
rect 379514 326408 379520 326460
rect 379572 326448 379578 326460
rect 380526 326448 380532 326460
rect 379572 326420 380532 326448
rect 379572 326408 379578 326420
rect 380526 326408 380532 326420
rect 380584 326408 380590 326460
rect 380894 326408 380900 326460
rect 380952 326448 380958 326460
rect 381998 326448 382004 326460
rect 380952 326420 382004 326448
rect 380952 326408 380958 326420
rect 381998 326408 382004 326420
rect 382056 326408 382062 326460
rect 383746 326408 383752 326460
rect 383804 326448 383810 326460
rect 384574 326448 384580 326460
rect 383804 326420 384580 326448
rect 383804 326408 383810 326420
rect 384574 326408 384580 326420
rect 384632 326408 384638 326460
rect 385218 326408 385224 326460
rect 385276 326448 385282 326460
rect 385678 326448 385684 326460
rect 385276 326420 385684 326448
rect 385276 326408 385282 326420
rect 385678 326408 385684 326420
rect 385736 326408 385742 326460
rect 386598 326408 386604 326460
rect 386656 326448 386662 326460
rect 387518 326448 387524 326460
rect 386656 326420 387524 326448
rect 386656 326408 386662 326420
rect 387518 326408 387524 326420
rect 387576 326408 387582 326460
rect 387886 326408 387892 326460
rect 387944 326448 387950 326460
rect 388254 326448 388260 326460
rect 387944 326420 388260 326448
rect 387944 326408 387950 326420
rect 388254 326408 388260 326420
rect 388312 326408 388318 326460
rect 401686 326408 401692 326460
rect 401744 326448 401750 326460
rect 402514 326448 402520 326460
rect 401744 326420 402520 326448
rect 401744 326408 401750 326420
rect 402514 326408 402520 326420
rect 402572 326408 402578 326460
rect 403066 326408 403072 326460
rect 403124 326448 403130 326460
rect 403526 326448 403532 326460
rect 403124 326420 403532 326448
rect 403124 326408 403130 326420
rect 403526 326408 403532 326420
rect 403584 326408 403590 326460
rect 404446 326408 404452 326460
rect 404504 326448 404510 326460
rect 404630 326448 404636 326460
rect 404504 326420 404636 326448
rect 404504 326408 404510 326420
rect 404630 326408 404636 326420
rect 404688 326408 404694 326460
rect 405918 326408 405924 326460
rect 405976 326448 405982 326460
rect 406470 326448 406476 326460
rect 405976 326420 406476 326448
rect 405976 326408 405982 326420
rect 406470 326408 406476 326420
rect 406528 326408 406534 326460
rect 407114 326408 407120 326460
rect 407172 326448 407178 326460
rect 407574 326448 407580 326460
rect 407172 326420 407580 326448
rect 407172 326408 407178 326420
rect 407574 326408 407580 326420
rect 407632 326408 407638 326460
rect 11698 326340 11704 326392
rect 11756 326380 11762 326392
rect 237006 326380 237012 326392
rect 11756 326352 237012 326380
rect 11756 326340 11762 326352
rect 237006 326340 237012 326352
rect 237064 326340 237070 326392
rect 237374 326340 237380 326392
rect 237432 326380 237438 326392
rect 238110 326380 238116 326392
rect 237432 326352 238116 326380
rect 237432 326340 237438 326352
rect 238110 326340 238116 326352
rect 238168 326340 238174 326392
rect 238754 326340 238760 326392
rect 238812 326380 238818 326392
rect 239582 326380 239588 326392
rect 238812 326352 239588 326380
rect 238812 326340 238818 326352
rect 239582 326340 239588 326352
rect 239640 326340 239646 326392
rect 240226 326340 240232 326392
rect 240284 326380 240290 326392
rect 240686 326380 240692 326392
rect 240284 326352 240692 326380
rect 240284 326340 240290 326352
rect 240686 326340 240692 326352
rect 240744 326340 240750 326392
rect 241606 326340 241612 326392
rect 241664 326380 241670 326392
rect 242158 326380 242164 326392
rect 241664 326352 242164 326380
rect 241664 326340 241670 326352
rect 242158 326340 242164 326352
rect 242216 326340 242222 326392
rect 274634 326340 274640 326392
rect 274692 326380 274698 326392
rect 275002 326380 275008 326392
rect 274692 326352 275008 326380
rect 274692 326340 274698 326352
rect 275002 326340 275008 326352
rect 275060 326340 275066 326392
rect 276014 326340 276020 326392
rect 276072 326380 276078 326392
rect 276474 326380 276480 326392
rect 276072 326352 276480 326380
rect 276072 326340 276078 326352
rect 276474 326340 276480 326352
rect 276532 326340 276538 326392
rect 277486 326340 277492 326392
rect 277544 326380 277550 326392
rect 278314 326380 278320 326392
rect 277544 326352 278320 326380
rect 277544 326340 277550 326352
rect 278314 326340 278320 326352
rect 278372 326340 278378 326392
rect 278958 326340 278964 326392
rect 279016 326380 279022 326392
rect 279418 326380 279424 326392
rect 279016 326352 279424 326380
rect 279016 326340 279022 326352
rect 279418 326340 279424 326352
rect 279476 326340 279482 326392
rect 280338 326340 280344 326392
rect 280396 326380 280402 326392
rect 281258 326380 281264 326392
rect 280396 326352 281264 326380
rect 280396 326340 280402 326352
rect 281258 326340 281264 326352
rect 281316 326340 281322 326392
rect 281534 326340 281540 326392
rect 281592 326380 281598 326392
rect 281994 326380 282000 326392
rect 281592 326352 282000 326380
rect 281592 326340 281598 326352
rect 281994 326340 282000 326352
rect 282052 326340 282058 326392
rect 304994 326340 305000 326392
rect 305052 326380 305058 326392
rect 306098 326380 306104 326392
rect 305052 326352 306104 326380
rect 305052 326340 305058 326352
rect 306098 326340 306104 326352
rect 306156 326340 306162 326392
rect 306558 326340 306564 326392
rect 306616 326380 306622 326392
rect 307478 326380 307484 326392
rect 306616 326352 307484 326380
rect 306616 326340 306622 326352
rect 307478 326340 307484 326352
rect 307536 326340 307542 326392
rect 309318 326340 309324 326392
rect 309376 326380 309382 326392
rect 310054 326380 310060 326392
rect 309376 326352 310060 326380
rect 309376 326340 309382 326352
rect 310054 326340 310060 326352
rect 310112 326340 310118 326392
rect 310606 326340 310612 326392
rect 310664 326380 310670 326392
rect 311158 326380 311164 326392
rect 310664 326352 311164 326380
rect 310664 326340 310670 326352
rect 311158 326340 311164 326352
rect 311216 326340 311222 326392
rect 321554 326340 321560 326392
rect 321612 326380 321618 326392
rect 322474 326380 322480 326392
rect 321612 326352 322480 326380
rect 321612 326340 321618 326352
rect 322474 326340 322480 326352
rect 322532 326340 322538 326392
rect 322934 326340 322940 326392
rect 322992 326380 322998 326392
rect 323578 326380 323584 326392
rect 322992 326352 323584 326380
rect 322992 326340 322998 326352
rect 323578 326340 323584 326352
rect 323636 326340 323642 326392
rect 327074 326340 327080 326392
rect 327132 326380 327138 326392
rect 327994 326380 328000 326392
rect 327132 326352 328000 326380
rect 327132 326340 327138 326352
rect 327994 326340 328000 326352
rect 328052 326340 328058 326392
rect 328638 326340 328644 326392
rect 328696 326380 328702 326392
rect 329466 326380 329472 326392
rect 328696 326352 329472 326380
rect 328696 326340 328702 326352
rect 329466 326340 329472 326352
rect 329524 326340 329530 326392
rect 329834 326340 329840 326392
rect 329892 326380 329898 326392
rect 330202 326380 330208 326392
rect 329892 326352 330208 326380
rect 329892 326340 329898 326352
rect 330202 326340 330208 326352
rect 330260 326340 330266 326392
rect 340966 326340 340972 326392
rect 341024 326380 341030 326392
rect 341886 326380 341892 326392
rect 341024 326352 341892 326380
rect 341024 326340 341030 326352
rect 341886 326340 341892 326352
rect 341944 326340 341950 326392
rect 342346 326340 342352 326392
rect 342404 326380 342410 326392
rect 343266 326380 343272 326392
rect 342404 326352 343272 326380
rect 342404 326340 342410 326352
rect 343266 326340 343272 326352
rect 343324 326340 343330 326392
rect 346486 326340 346492 326392
rect 346544 326380 346550 326392
rect 347406 326380 347412 326392
rect 346544 326352 347412 326380
rect 346544 326340 346550 326352
rect 347406 326340 347412 326352
rect 347464 326340 347470 326392
rect 350534 326340 350540 326392
rect 350592 326380 350598 326392
rect 351362 326380 351368 326392
rect 350592 326352 351368 326380
rect 350592 326340 350598 326352
rect 351362 326340 351368 326352
rect 351420 326340 351426 326392
rect 354766 326340 354772 326392
rect 354824 326380 354830 326392
rect 355318 326380 355324 326392
rect 354824 326352 355324 326380
rect 354824 326340 354830 326352
rect 355318 326340 355324 326352
rect 355376 326340 355382 326392
rect 356054 326340 356060 326392
rect 356112 326380 356118 326392
rect 357158 326380 357164 326392
rect 356112 326352 357164 326380
rect 356112 326340 356118 326352
rect 357158 326340 357164 326352
rect 357216 326340 357222 326392
rect 357526 326340 357532 326392
rect 357584 326380 357590 326392
rect 358262 326380 358268 326392
rect 357584 326352 358268 326380
rect 357584 326340 357590 326352
rect 358262 326340 358268 326352
rect 358320 326340 358326 326392
rect 364610 326340 364616 326392
rect 364668 326380 364674 326392
rect 419534 326380 419540 326392
rect 364668 326352 419540 326380
rect 364668 326340 364674 326352
rect 419534 326340 419540 326352
rect 419592 326340 419598 326392
rect 241514 326272 241520 326324
rect 241572 326312 241578 326324
rect 242526 326312 242532 326324
rect 241572 326284 242532 326312
rect 241572 326272 241578 326284
rect 242526 326272 242532 326284
rect 242584 326272 242590 326324
rect 278774 326272 278780 326324
rect 278832 326312 278838 326324
rect 279786 326312 279792 326324
rect 278832 326284 279792 326312
rect 278832 326272 278838 326284
rect 279786 326272 279792 326284
rect 279844 326272 279850 326324
rect 280154 326272 280160 326324
rect 280212 326312 280218 326324
rect 280890 326312 280896 326324
rect 280212 326284 280896 326312
rect 280212 326272 280218 326284
rect 280890 326272 280896 326284
rect 280948 326272 280954 326324
rect 371234 326272 371240 326324
rect 371292 326312 371298 326324
rect 371786 326312 371792 326324
rect 371292 326284 371792 326312
rect 371292 326272 371298 326284
rect 371786 326272 371792 326284
rect 371844 326272 371850 326324
rect 378226 326272 378232 326324
rect 378284 326312 378290 326324
rect 379146 326312 379152 326324
rect 378284 326284 379152 326312
rect 378284 326272 378290 326284
rect 379146 326272 379152 326284
rect 379204 326272 379210 326324
rect 387794 326272 387800 326324
rect 387852 326312 387858 326324
rect 388622 326312 388628 326324
rect 387852 326284 388628 326312
rect 387852 326272 387858 326284
rect 388622 326272 388628 326284
rect 388680 326272 388686 326324
rect 402974 326272 402980 326324
rect 403032 326312 403038 326324
rect 403894 326312 403900 326324
rect 403032 326284 403900 326312
rect 403032 326272 403038 326284
rect 403894 326272 403900 326284
rect 403952 326272 403958 326324
rect 405734 326272 405740 326324
rect 405792 326312 405798 326324
rect 406838 326312 406844 326324
rect 405792 326284 406844 326312
rect 405792 326272 405798 326284
rect 406838 326272 406844 326284
rect 406896 326272 406902 326324
rect 407206 326272 407212 326324
rect 407264 326312 407270 326324
rect 407942 326312 407948 326324
rect 407264 326284 407948 326312
rect 407264 326272 407270 326284
rect 407942 326272 407948 326284
rect 408000 326272 408006 326324
rect 242894 326000 242900 326052
rect 242952 326040 242958 326052
rect 243630 326040 243636 326052
rect 242952 326012 243636 326040
rect 242952 326000 242958 326012
rect 243630 326000 243636 326012
rect 243688 326000 243694 326052
rect 176654 324980 176660 325032
rect 176712 325020 176718 325032
rect 289906 325020 289912 325032
rect 176712 324992 289912 325020
rect 176712 324980 176718 324992
rect 289906 324980 289912 324992
rect 289964 324980 289970 325032
rect 160094 324912 160100 324964
rect 160152 324952 160158 324964
rect 276750 324952 276756 324964
rect 160152 324924 276756 324952
rect 160152 324912 160158 324924
rect 276750 324912 276756 324924
rect 276808 324912 276814 324964
rect 365990 324912 365996 324964
rect 366048 324952 366054 324964
rect 423674 324952 423680 324964
rect 366048 324924 423680 324952
rect 366048 324912 366054 324924
rect 423674 324912 423680 324924
rect 423732 324912 423738 324964
rect 292574 324844 292580 324896
rect 292632 324884 292638 324896
rect 292758 324884 292764 324896
rect 292632 324856 292764 324884
rect 292632 324844 292638 324856
rect 292758 324844 292764 324856
rect 292816 324844 292822 324896
rect 347774 323824 347780 323876
rect 347832 323864 347838 323876
rect 348786 323864 348792 323876
rect 347832 323836 348792 323864
rect 347832 323824 347838 323836
rect 348786 323824 348792 323836
rect 348844 323824 348850 323876
rect 386506 323824 386512 323876
rect 386564 323864 386570 323876
rect 387150 323864 387156 323876
rect 386564 323836 387156 323864
rect 386564 323824 386570 323836
rect 387150 323824 387156 323836
rect 387208 323824 387214 323876
rect 385034 323688 385040 323740
rect 385092 323728 385098 323740
rect 386046 323728 386052 323740
rect 385092 323700 386052 323728
rect 385092 323688 385098 323700
rect 386046 323688 386052 323700
rect 386104 323688 386110 323740
rect 128354 323620 128360 323672
rect 128412 323660 128418 323672
rect 274818 323660 274824 323672
rect 128412 323632 274824 323660
rect 128412 323620 128418 323632
rect 274818 323620 274824 323632
rect 274876 323620 274882 323672
rect 26234 323552 26240 323604
rect 26292 323592 26298 323604
rect 243170 323592 243176 323604
rect 26292 323564 243176 323592
rect 26292 323552 26298 323564
rect 243170 323552 243176 323564
rect 243228 323552 243234 323604
rect 305178 323552 305184 323604
rect 305236 323592 305242 323604
rect 305362 323592 305368 323604
rect 305236 323564 305368 323592
rect 305236 323552 305242 323564
rect 305362 323552 305368 323564
rect 305420 323552 305426 323604
rect 358814 323552 358820 323604
rect 358872 323592 358878 323604
rect 359090 323592 359096 323604
rect 358872 323564 359096 323592
rect 358872 323552 358878 323564
rect 359090 323552 359096 323564
rect 359148 323552 359154 323604
rect 378134 323552 378140 323604
rect 378192 323592 378198 323604
rect 378410 323592 378416 323604
rect 378192 323564 378416 323592
rect 378192 323552 378198 323564
rect 378410 323552 378416 323564
rect 378468 323552 378474 323604
rect 398466 323552 398472 323604
rect 398524 323592 398530 323604
rect 529934 323592 529940 323604
rect 398524 323564 529940 323592
rect 398524 323552 398530 323564
rect 529934 323552 529940 323564
rect 529992 323552 529998 323604
rect 302418 323280 302424 323332
rect 302476 323320 302482 323332
rect 303154 323320 303160 323332
rect 302476 323292 303160 323320
rect 302476 323280 302482 323292
rect 303154 323280 303160 323292
rect 303212 323280 303218 323332
rect 343634 323280 343640 323332
rect 343692 323320 343698 323332
rect 344370 323320 344376 323332
rect 343692 323292 344376 323320
rect 343692 323280 343698 323292
rect 344370 323280 344376 323292
rect 344428 323280 344434 323332
rect 358906 323212 358912 323264
rect 358964 323252 358970 323264
rect 359734 323252 359740 323264
rect 358964 323224 359740 323252
rect 358964 323212 358970 323224
rect 359734 323212 359740 323224
rect 359792 323212 359798 323264
rect 305086 322464 305092 322516
rect 305144 322504 305150 322516
rect 305730 322504 305736 322516
rect 305144 322476 305736 322504
rect 305144 322464 305150 322476
rect 305730 322464 305736 322476
rect 305788 322464 305794 322516
rect 403158 322464 403164 322516
rect 403216 322504 403222 322516
rect 403342 322504 403348 322516
rect 403216 322476 403348 322504
rect 403216 322464 403222 322476
rect 403342 322464 403348 322476
rect 403400 322464 403406 322516
rect 189074 322260 189080 322312
rect 189132 322300 189138 322312
rect 291930 322300 291936 322312
rect 189132 322272 291936 322300
rect 189132 322260 189138 322272
rect 291930 322260 291936 322272
rect 291988 322260 291994 322312
rect 51074 322192 51080 322244
rect 51132 322232 51138 322244
rect 250530 322232 250536 322244
rect 51132 322204 250536 322232
rect 51132 322192 51138 322204
rect 250530 322192 250536 322204
rect 250588 322192 250594 322244
rect 345014 322192 345020 322244
rect 345072 322232 345078 322244
rect 345842 322232 345848 322244
rect 345072 322204 345848 322232
rect 345072 322192 345078 322204
rect 345842 322192 345848 322204
rect 345900 322192 345906 322244
rect 398926 322192 398932 322244
rect 398984 322232 398990 322244
rect 532694 322232 532700 322244
rect 398984 322204 532700 322232
rect 398984 322192 398990 322204
rect 532694 322192 532700 322204
rect 532752 322192 532758 322244
rect 273346 322056 273352 322108
rect 273404 322096 273410 322108
rect 273898 322096 273904 322108
rect 273404 322068 273904 322096
rect 273404 322056 273410 322068
rect 273898 322056 273904 322068
rect 273956 322056 273962 322108
rect 347866 321512 347872 321564
rect 347924 321552 347930 321564
rect 348050 321552 348056 321564
rect 347924 321524 348056 321552
rect 347924 321512 347930 321524
rect 348050 321512 348056 321524
rect 348108 321512 348114 321564
rect 367370 320900 367376 320952
rect 367428 320940 367434 320952
rect 427814 320940 427820 320952
rect 367428 320912 427820 320940
rect 367428 320900 367434 320912
rect 427814 320900 427820 320912
rect 427872 320900 427878 320952
rect 215294 320832 215300 320884
rect 215352 320872 215358 320884
rect 301314 320872 301320 320884
rect 215352 320844 301320 320872
rect 215352 320832 215358 320844
rect 301314 320832 301320 320844
rect 301372 320832 301378 320884
rect 385310 320832 385316 320884
rect 385368 320872 385374 320884
rect 487154 320872 487160 320884
rect 385368 320844 487160 320872
rect 385368 320832 385374 320844
rect 487154 320832 487160 320844
rect 487212 320832 487218 320884
rect 248414 320764 248420 320816
rect 248472 320804 248478 320816
rect 248598 320804 248604 320816
rect 248472 320776 248604 320804
rect 248472 320764 248478 320776
rect 248598 320764 248604 320776
rect 248656 320764 248662 320816
rect 3510 320084 3516 320136
rect 3568 320124 3574 320136
rect 232498 320124 232504 320136
rect 3568 320096 232504 320124
rect 3568 320084 3574 320096
rect 232498 320084 232504 320096
rect 232556 320084 232562 320136
rect 325786 319472 325792 319524
rect 325844 319512 325850 319524
rect 325970 319512 325976 319524
rect 325844 319484 325976 319512
rect 325844 319472 325850 319484
rect 325970 319472 325976 319484
rect 326028 319472 326034 319524
rect 369210 319472 369216 319524
rect 369268 319512 369274 319524
rect 434714 319512 434720 319524
rect 369268 319484 434720 319512
rect 369268 319472 369274 319484
rect 434714 319472 434720 319484
rect 434772 319472 434778 319524
rect 205634 319404 205640 319456
rect 205692 319444 205698 319456
rect 298278 319444 298284 319456
rect 205692 319416 298284 319444
rect 205692 319404 205698 319416
rect 298278 319404 298284 319416
rect 298336 319404 298342 319456
rect 386690 319404 386696 319456
rect 386748 319444 386754 319456
rect 489914 319444 489920 319456
rect 386748 319416 489920 319444
rect 386748 319404 386754 319416
rect 489914 319404 489920 319416
rect 489972 319404 489978 319456
rect 371510 318112 371516 318164
rect 371568 318152 371574 318164
rect 441614 318152 441620 318164
rect 371568 318124 441620 318152
rect 371568 318112 371574 318124
rect 441614 318112 441620 318124
rect 441672 318112 441678 318164
rect 219434 318044 219440 318096
rect 219492 318084 219498 318096
rect 302326 318084 302332 318096
rect 219492 318056 302332 318084
rect 219492 318044 219498 318056
rect 302326 318044 302332 318056
rect 302384 318044 302390 318096
rect 386598 318044 386604 318096
rect 386656 318084 386662 318096
rect 494054 318084 494060 318096
rect 386656 318056 494060 318084
rect 386656 318044 386662 318056
rect 494054 318044 494060 318056
rect 494112 318044 494118 318096
rect 223574 316684 223580 316736
rect 223632 316724 223638 316736
rect 303798 316724 303804 316736
rect 223632 316696 303804 316724
rect 223632 316684 223638 316696
rect 303798 316684 303804 316696
rect 303856 316684 303862 316736
rect 387794 316684 387800 316736
rect 387852 316724 387858 316736
rect 498194 316724 498200 316736
rect 387852 316696 498200 316724
rect 387852 316684 387858 316696
rect 498194 316684 498200 316696
rect 498252 316684 498258 316736
rect 226334 315256 226340 315308
rect 226392 315296 226398 315308
rect 305270 315296 305276 315308
rect 226392 315268 305276 315296
rect 226392 315256 226398 315268
rect 305270 315256 305276 315268
rect 305328 315256 305334 315308
rect 394694 315256 394700 315308
rect 394752 315296 394758 315308
rect 518894 315296 518900 315308
rect 394752 315268 518900 315296
rect 394752 315256 394758 315268
rect 518894 315256 518900 315268
rect 518952 315256 518958 315308
rect 118694 313896 118700 313948
rect 118752 313936 118758 313948
rect 272058 313936 272064 313948
rect 118752 313908 272064 313936
rect 118752 313896 118758 313908
rect 272058 313896 272064 313908
rect 272116 313896 272122 313948
rect 391934 313896 391940 313948
rect 391992 313936 391998 313948
rect 511994 313936 512000 313948
rect 391992 313908 512000 313936
rect 391992 313896 391998 313908
rect 511994 313896 512000 313908
rect 512052 313896 512058 313948
rect 171134 312604 171140 312656
rect 171192 312644 171198 312656
rect 286410 312644 286416 312656
rect 171192 312616 286416 312644
rect 171192 312604 171198 312616
rect 286410 312604 286416 312616
rect 286468 312604 286474 312656
rect 69014 312536 69020 312588
rect 69072 312576 69078 312588
rect 255590 312576 255596 312588
rect 69072 312548 255596 312576
rect 69072 312536 69078 312548
rect 255590 312536 255596 312548
rect 255648 312536 255654 312588
rect 370038 312536 370044 312588
rect 370096 312576 370102 312588
rect 438854 312576 438860 312588
rect 370096 312548 438860 312576
rect 370096 312536 370102 312548
rect 438854 312536 438860 312548
rect 438912 312536 438918 312588
rect 122834 311108 122840 311160
rect 122892 311148 122898 311160
rect 271966 311148 271972 311160
rect 122892 311120 271972 311148
rect 122892 311108 122898 311120
rect 271966 311108 271972 311120
rect 272024 311108 272030 311160
rect 400306 311108 400312 311160
rect 400364 311148 400370 311160
rect 536834 311148 536840 311160
rect 400364 311120 536840 311148
rect 400364 311108 400370 311120
rect 536834 311108 536840 311120
rect 536892 311108 536898 311160
rect 135254 309748 135260 309800
rect 135312 309788 135318 309800
rect 276198 309788 276204 309800
rect 135312 309760 276204 309788
rect 135312 309748 135318 309760
rect 276198 309748 276204 309760
rect 276256 309748 276262 309800
rect 406010 309748 406016 309800
rect 406068 309788 406074 309800
rect 554774 309788 554780 309800
rect 406068 309760 554780 309788
rect 406068 309748 406074 309760
rect 554774 309748 554780 309760
rect 554832 309748 554838 309800
rect 132494 308456 132500 308508
rect 132552 308496 132558 308508
rect 274818 308496 274824 308508
rect 132552 308468 274824 308496
rect 132552 308456 132558 308468
rect 274818 308456 274824 308468
rect 274876 308456 274882 308508
rect 74534 308388 74540 308440
rect 74592 308428 74598 308440
rect 258350 308428 258356 308440
rect 74592 308400 258356 308428
rect 74592 308388 74598 308400
rect 258350 308388 258356 308400
rect 258408 308388 258414 308440
rect 408678 308388 408684 308440
rect 408736 308428 408742 308440
rect 564434 308428 564440 308440
rect 408736 308400 564440 308428
rect 408736 308388 408742 308400
rect 564434 308388 564440 308400
rect 564492 308388 564498 308440
rect 207014 307096 207020 307148
rect 207072 307136 207078 307148
rect 294598 307136 294604 307148
rect 207072 307108 294604 307136
rect 207072 307096 207078 307108
rect 294598 307096 294604 307108
rect 294656 307096 294662 307148
rect 64874 307028 64880 307080
rect 64932 307068 64938 307080
rect 254026 307068 254032 307080
rect 64932 307040 254032 307068
rect 64932 307028 64938 307040
rect 254026 307028 254032 307040
rect 254084 307028 254090 307080
rect 381078 307028 381084 307080
rect 381136 307068 381142 307080
rect 473354 307068 473360 307080
rect 381136 307040 473360 307068
rect 381136 307028 381142 307040
rect 473354 307028 473360 307040
rect 473412 307028 473418 307080
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 383010 306320 383016 306332
rect 3384 306292 383016 306320
rect 3384 306280 3390 306292
rect 383010 306280 383016 306292
rect 383068 306280 383074 306332
rect 379606 305668 379612 305720
rect 379664 305708 379670 305720
rect 470594 305708 470600 305720
rect 379664 305680 470600 305708
rect 379664 305668 379670 305680
rect 470594 305668 470600 305680
rect 470652 305668 470658 305720
rect 390830 305600 390836 305652
rect 390888 305640 390894 305652
rect 505094 305640 505100 305652
rect 390888 305612 505100 305640
rect 390888 305600 390894 305612
rect 505094 305600 505100 305612
rect 505152 305600 505158 305652
rect 209774 304308 209780 304360
rect 209832 304348 209838 304360
rect 297450 304348 297456 304360
rect 209832 304320 297456 304348
rect 209832 304308 209838 304320
rect 297450 304308 297456 304320
rect 297508 304308 297514 304360
rect 53834 304240 53840 304292
rect 53892 304280 53898 304292
rect 251358 304280 251364 304292
rect 53892 304252 251364 304280
rect 53892 304240 53898 304252
rect 251358 304240 251364 304252
rect 251416 304240 251422 304292
rect 413278 304240 413284 304292
rect 413336 304280 413342 304292
rect 572806 304280 572812 304292
rect 413336 304252 572812 304280
rect 413336 304240 413342 304252
rect 572806 304240 572812 304252
rect 572864 304240 572870 304292
rect 179414 302948 179420 303000
rect 179472 302988 179478 303000
rect 287698 302988 287704 303000
rect 179472 302960 287704 302988
rect 179472 302948 179478 302960
rect 287698 302948 287704 302960
rect 287756 302948 287762 303000
rect 15838 302880 15844 302932
rect 15896 302920 15902 302932
rect 237650 302920 237656 302932
rect 15896 302892 237656 302920
rect 15896 302880 15902 302892
rect 237650 302880 237656 302892
rect 237708 302880 237714 302932
rect 146294 301452 146300 301504
rect 146352 301492 146358 301504
rect 280430 301492 280436 301504
rect 146352 301464 280436 301492
rect 146352 301452 146358 301464
rect 280430 301452 280436 301464
rect 280488 301452 280494 301504
rect 393498 301452 393504 301504
rect 393556 301492 393562 301504
rect 513374 301492 513380 301504
rect 393556 301464 513380 301492
rect 393556 301452 393562 301464
rect 513374 301452 513380 301464
rect 513432 301452 513438 301504
rect 143534 300092 143540 300144
rect 143592 300132 143598 300144
rect 279050 300132 279056 300144
rect 143592 300104 279056 300132
rect 143592 300092 143598 300104
rect 279050 300092 279056 300104
rect 279108 300092 279114 300144
rect 397546 300092 397552 300144
rect 397604 300132 397610 300144
rect 527174 300132 527180 300144
rect 397604 300104 527180 300132
rect 397604 300092 397610 300104
rect 527174 300092 527180 300104
rect 527232 300092 527238 300144
rect 424410 299412 424416 299464
rect 424468 299452 424474 299464
rect 580166 299452 580172 299464
rect 424468 299424 580172 299452
rect 424468 299412 424474 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 361666 298732 361672 298784
rect 361724 298772 361730 298784
rect 409874 298772 409880 298784
rect 361724 298744 409880 298772
rect 361724 298732 361730 298744
rect 409874 298732 409880 298744
rect 409932 298732 409938 298784
rect 403250 297372 403256 297424
rect 403308 297412 403314 297424
rect 543734 297412 543740 297424
rect 403308 297384 543740 297412
rect 403308 297372 403314 297384
rect 543734 297372 543740 297384
rect 543792 297372 543798 297424
rect 402974 295944 402980 295996
rect 403032 295984 403038 295996
rect 547874 295984 547880 295996
rect 403032 295956 547880 295984
rect 403032 295944 403038 295956
rect 547874 295944 547880 295956
rect 547932 295944 547938 295996
rect 407298 294584 407304 294636
rect 407356 294624 407362 294636
rect 557534 294624 557540 294636
rect 407356 294596 557540 294624
rect 407356 294584 407362 294596
rect 557534 294584 557540 294596
rect 557592 294584 557598 294636
rect 2866 293904 2872 293956
rect 2924 293944 2930 293956
rect 18598 293944 18604 293956
rect 2924 293916 18604 293944
rect 2924 293904 2930 293916
rect 18598 293904 18604 293916
rect 18656 293904 18662 293956
rect 410150 293224 410156 293276
rect 410208 293264 410214 293276
rect 568574 293264 568580 293276
rect 410208 293236 568580 293264
rect 410208 293224 410214 293236
rect 568574 293224 568580 293236
rect 568632 293224 568638 293276
rect 154574 291796 154580 291848
rect 154632 291836 154638 291848
rect 283190 291836 283196 291848
rect 154632 291808 283196 291836
rect 154632 291796 154638 291808
rect 283190 291796 283196 291808
rect 283248 291796 283254 291848
rect 408586 291796 408592 291848
rect 408644 291836 408650 291848
rect 563054 291836 563060 291848
rect 408644 291808 563060 291836
rect 408644 291796 408650 291808
rect 563054 291796 563060 291808
rect 563112 291796 563118 291848
rect 136634 290436 136640 290488
rect 136692 290476 136698 290488
rect 277578 290476 277584 290488
rect 136692 290448 277584 290476
rect 136692 290436 136698 290448
rect 277578 290436 277584 290448
rect 277636 290436 277642 290488
rect 410058 290436 410064 290488
rect 410116 290476 410122 290488
rect 565814 290476 565820 290488
rect 410116 290448 565820 290476
rect 410116 290436 410122 290448
rect 565814 290436 565820 290448
rect 565872 290436 565878 290488
rect 157334 289144 157340 289196
rect 157392 289184 157398 289196
rect 283098 289184 283104 289196
rect 157392 289156 283104 289184
rect 157392 289144 157398 289156
rect 283098 289144 283104 289156
rect 283156 289144 283162 289196
rect 81434 289076 81440 289128
rect 81492 289116 81498 289128
rect 259730 289116 259736 289128
rect 81492 289088 259736 289116
rect 81492 289076 81498 289088
rect 259730 289076 259736 289088
rect 259788 289076 259794 289128
rect 411438 289076 411444 289128
rect 411496 289116 411502 289128
rect 571978 289116 571984 289128
rect 411496 289088 571984 289116
rect 411496 289076 411502 289088
rect 571978 289076 571984 289088
rect 572036 289076 572042 289128
rect 139394 287648 139400 287700
rect 139452 287688 139458 287700
rect 276658 287688 276664 287700
rect 139452 287660 276664 287688
rect 139452 287648 139458 287660
rect 276658 287648 276664 287660
rect 276716 287648 276722 287700
rect 397454 287648 397460 287700
rect 397512 287688 397518 287700
rect 528554 287688 528560 287700
rect 397512 287660 528560 287688
rect 397512 287648 397518 287660
rect 528554 287648 528560 287660
rect 528612 287648 528618 287700
rect 178034 286356 178040 286408
rect 178092 286396 178098 286408
rect 289170 286396 289176 286408
rect 178092 286368 289176 286396
rect 178092 286356 178098 286368
rect 289170 286356 289176 286368
rect 289228 286356 289234 286408
rect 354950 286356 354956 286408
rect 355008 286396 355014 286408
rect 387794 286396 387800 286408
rect 355008 286368 387800 286396
rect 355008 286356 355014 286368
rect 387794 286356 387800 286368
rect 387852 286356 387858 286408
rect 6270 286288 6276 286340
rect 6328 286328 6334 286340
rect 236086 286328 236092 286340
rect 6328 286300 236092 286328
rect 6328 286288 6334 286300
rect 236086 286288 236092 286300
rect 236144 286288 236150 286340
rect 376938 286288 376944 286340
rect 376996 286328 377002 286340
rect 462314 286328 462320 286340
rect 376996 286300 462320 286328
rect 376996 286288 377002 286300
rect 462314 286288 462320 286300
rect 462372 286288 462378 286340
rect 182174 284996 182180 285048
rect 182232 285036 182238 285048
rect 286318 285036 286324 285048
rect 182232 285008 286324 285036
rect 182232 284996 182238 285008
rect 286318 284996 286324 285008
rect 286376 284996 286382 285048
rect 356330 284996 356336 285048
rect 356388 285036 356394 285048
rect 394694 285036 394700 285048
rect 356388 285008 394700 285036
rect 356388 284996 356394 285008
rect 394694 284996 394700 285008
rect 394752 284996 394758 285048
rect 40034 284928 40040 284980
rect 40092 284968 40098 284980
rect 246298 284968 246304 284980
rect 40092 284940 246304 284968
rect 40092 284928 40098 284940
rect 246298 284928 246304 284940
rect 246356 284928 246362 284980
rect 285674 284928 285680 284980
rect 285732 284968 285738 284980
rect 323210 284968 323216 284980
rect 285732 284940 323216 284968
rect 285732 284928 285738 284940
rect 323210 284928 323216 284940
rect 323268 284928 323274 284980
rect 378410 284928 378416 284980
rect 378468 284968 378474 284980
rect 465166 284968 465172 284980
rect 378468 284940 465172 284968
rect 378468 284928 378474 284940
rect 465166 284928 465172 284940
rect 465224 284928 465230 284980
rect 184934 283636 184940 283688
rect 184992 283676 184998 283688
rect 291378 283676 291384 283688
rect 184992 283648 291384 283676
rect 184992 283636 184998 283648
rect 291378 283636 291384 283648
rect 291436 283636 291442 283688
rect 360470 283636 360476 283688
rect 360528 283676 360534 283688
rect 408586 283676 408592 283688
rect 360528 283648 408592 283676
rect 360528 283636 360534 283648
rect 408586 283636 408592 283648
rect 408644 283636 408650 283688
rect 35894 283568 35900 283620
rect 35952 283608 35958 283620
rect 244918 283608 244924 283620
rect 35952 283580 244924 283608
rect 35952 283568 35958 283580
rect 244918 283568 244924 283580
rect 244976 283568 244982 283620
rect 390738 283568 390744 283620
rect 390796 283608 390802 283620
rect 506474 283608 506480 283620
rect 390796 283580 506480 283608
rect 390796 283568 390802 283580
rect 506474 283568 506480 283580
rect 506532 283568 506538 283620
rect 195974 282208 195980 282260
rect 196032 282248 196038 282260
rect 295518 282248 295524 282260
rect 196032 282220 295524 282248
rect 196032 282208 196038 282220
rect 295518 282208 295524 282220
rect 295576 282208 295582 282260
rect 363230 282208 363236 282260
rect 363288 282248 363294 282260
rect 415394 282248 415400 282260
rect 363288 282220 415400 282248
rect 363288 282208 363294 282220
rect 415394 282208 415400 282220
rect 415452 282208 415458 282260
rect 20714 282140 20720 282192
rect 20772 282180 20778 282192
rect 241790 282180 241796 282192
rect 20772 282152 241796 282180
rect 20772 282140 20778 282152
rect 241790 282140 241796 282152
rect 241848 282140 241854 282192
rect 394878 282140 394884 282192
rect 394936 282180 394942 282192
rect 520274 282180 520280 282192
rect 394936 282152 520280 282180
rect 394936 282140 394942 282152
rect 520274 282140 520280 282152
rect 520332 282140 520338 282192
rect 200114 280848 200120 280900
rect 200172 280888 200178 280900
rect 295978 280888 295984 280900
rect 200172 280860 295984 280888
rect 200172 280848 200178 280860
rect 295978 280848 295984 280860
rect 296036 280848 296042 280900
rect 365898 280848 365904 280900
rect 365956 280888 365962 280900
rect 423766 280888 423772 280900
rect 365956 280860 423772 280888
rect 365956 280848 365962 280860
rect 423766 280848 423772 280860
rect 423824 280848 423830 280900
rect 121454 280780 121460 280832
rect 121512 280820 121518 280832
rect 271138 280820 271144 280832
rect 121512 280792 271144 280820
rect 121512 280780 121518 280792
rect 271138 280780 271144 280792
rect 271196 280780 271202 280832
rect 404538 280780 404544 280832
rect 404596 280820 404602 280832
rect 552014 280820 552020 280832
rect 404596 280792 552020 280820
rect 404596 280780 404602 280792
rect 552014 280780 552020 280792
rect 552072 280780 552078 280832
rect 296714 279624 296720 279676
rect 296772 279664 296778 279676
rect 320818 279664 320824 279676
rect 296772 279636 320824 279664
rect 296772 279624 296778 279636
rect 320818 279624 320824 279636
rect 320876 279624 320882 279676
rect 202874 279488 202880 279540
rect 202932 279528 202938 279540
rect 296990 279528 296996 279540
rect 202932 279500 296996 279528
rect 202932 279488 202938 279500
rect 296990 279488 296996 279500
rect 297048 279488 297054 279540
rect 365806 279488 365812 279540
rect 365864 279528 365870 279540
rect 426434 279528 426440 279540
rect 365864 279500 426440 279528
rect 365864 279488 365870 279500
rect 426434 279488 426440 279500
rect 426492 279488 426498 279540
rect 96614 279420 96620 279472
rect 96672 279460 96678 279472
rect 264238 279460 264244 279472
rect 96672 279432 264244 279460
rect 96672 279420 96678 279432
rect 264238 279420 264244 279432
rect 264296 279420 264302 279472
rect 405918 279420 405924 279472
rect 405976 279460 405982 279472
rect 556154 279460 556160 279472
rect 405976 279432 556160 279460
rect 405976 279420 405982 279432
rect 556154 279420 556160 279432
rect 556212 279420 556218 279472
rect 213914 278060 213920 278112
rect 213972 278100 213978 278112
rect 300946 278100 300952 278112
rect 213972 278072 300952 278100
rect 213972 278060 213978 278072
rect 300946 278060 300952 278072
rect 301004 278060 301010 278112
rect 372798 278060 372804 278112
rect 372856 278100 372862 278112
rect 448514 278100 448520 278112
rect 372856 278072 448520 278100
rect 372856 278060 372862 278072
rect 448514 278060 448520 278072
rect 448572 278060 448578 278112
rect 89714 277992 89720 278044
rect 89772 278032 89778 278044
rect 262490 278032 262496 278044
rect 89772 278004 262496 278032
rect 89772 277992 89778 278004
rect 262490 277992 262496 278004
rect 262548 277992 262554 278044
rect 412818 277992 412824 278044
rect 412876 278032 412882 278044
rect 576118 278032 576124 278044
rect 412876 278004 576124 278032
rect 412876 277992 412882 278004
rect 576118 277992 576124 278004
rect 576176 277992 576182 278044
rect 220814 276700 220820 276752
rect 220872 276740 220878 276752
rect 302418 276740 302424 276752
rect 220872 276712 302424 276740
rect 220872 276700 220878 276712
rect 302418 276700 302424 276712
rect 302476 276700 302482 276752
rect 85574 276632 85580 276684
rect 85632 276672 85638 276684
rect 261110 276672 261116 276684
rect 85632 276644 261116 276672
rect 85632 276632 85638 276644
rect 261110 276632 261116 276644
rect 261168 276632 261174 276684
rect 374270 276632 374276 276684
rect 374328 276672 374334 276684
rect 451274 276672 451280 276684
rect 374328 276644 451280 276672
rect 374328 276632 374334 276644
rect 451274 276632 451280 276644
rect 451332 276632 451338 276684
rect 227714 275340 227720 275392
rect 227772 275380 227778 275392
rect 305178 275380 305184 275392
rect 227772 275352 305184 275380
rect 227772 275340 227778 275352
rect 305178 275340 305184 275352
rect 305236 275340 305242 275392
rect 4798 275272 4804 275324
rect 4856 275312 4862 275324
rect 234706 275312 234712 275324
rect 4856 275284 234712 275312
rect 4856 275272 4862 275284
rect 234706 275272 234712 275284
rect 234764 275272 234770 275324
rect 375558 275272 375564 275324
rect 375616 275312 375622 275324
rect 455414 275312 455420 275324
rect 375616 275284 455420 275312
rect 375616 275272 375622 275284
rect 455414 275272 455420 275284
rect 455472 275272 455478 275324
rect 274818 274048 274824 274100
rect 274876 274088 274882 274100
rect 319070 274088 319076 274100
rect 274876 274060 319076 274088
rect 274876 274048 274882 274060
rect 319070 274048 319076 274060
rect 319128 274048 319134 274100
rect 129734 273912 129740 273964
rect 129792 273952 129798 273964
rect 274634 273952 274640 273964
rect 129792 273924 274640 273952
rect 129792 273912 129798 273924
rect 274634 273912 274640 273924
rect 274692 273912 274698 273964
rect 376846 273912 376852 273964
rect 376904 273952 376910 273964
rect 458174 273952 458180 273964
rect 376904 273924 458180 273952
rect 376904 273912 376910 273924
rect 458174 273912 458180 273924
rect 458232 273912 458238 273964
rect 431218 273164 431224 273216
rect 431276 273204 431282 273216
rect 580166 273204 580172 273216
rect 431276 273176 580172 273204
rect 431276 273164 431282 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 150434 272484 150440 272536
rect 150492 272524 150498 272536
rect 280338 272524 280344 272536
rect 150492 272496 280344 272524
rect 150492 272484 150498 272496
rect 280338 272484 280344 272496
rect 280396 272484 280402 272536
rect 359090 272484 359096 272536
rect 359148 272524 359154 272536
rect 402974 272524 402980 272536
rect 359148 272496 402980 272524
rect 359148 272484 359154 272496
rect 402974 272484 402980 272496
rect 403032 272484 403038 272536
rect 153194 271124 153200 271176
rect 153252 271164 153258 271176
rect 281718 271164 281724 271176
rect 153252 271136 281724 271164
rect 153252 271124 153258 271136
rect 281718 271124 281724 271136
rect 281776 271124 281782 271176
rect 381538 271124 381544 271176
rect 381596 271164 381602 271176
rect 469214 271164 469220 271176
rect 381596 271136 469220 271164
rect 381596 271124 381602 271136
rect 469214 271124 469220 271136
rect 469272 271124 469278 271176
rect 161474 269764 161480 269816
rect 161532 269804 161538 269816
rect 284478 269804 284484 269816
rect 161532 269776 284484 269804
rect 161532 269764 161538 269776
rect 284478 269764 284484 269776
rect 284536 269764 284542 269816
rect 383838 269764 383844 269816
rect 383896 269804 383902 269816
rect 481634 269804 481640 269816
rect 383896 269776 481640 269804
rect 383896 269764 383902 269776
rect 481634 269764 481640 269776
rect 481692 269764 481698 269816
rect 165614 268336 165620 268388
rect 165672 268376 165678 268388
rect 285858 268376 285864 268388
rect 165672 268348 285864 268376
rect 165672 268336 165678 268348
rect 285858 268336 285864 268348
rect 285916 268336 285922 268388
rect 383746 268336 383752 268388
rect 383804 268376 383810 268388
rect 484394 268376 484400 268388
rect 383804 268348 484400 268376
rect 383804 268336 383810 268348
rect 484394 268336 484400 268348
rect 484452 268336 484458 268388
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 231210 267696 231216 267708
rect 3292 267668 231216 267696
rect 3292 267656 3298 267668
rect 231210 267656 231216 267668
rect 231268 267656 231274 267708
rect 222194 266976 222200 267028
rect 222252 267016 222258 267028
rect 303706 267016 303712 267028
rect 222252 266988 303712 267016
rect 222252 266976 222258 266988
rect 303706 266976 303712 266988
rect 303764 266976 303770 267028
rect 385218 266976 385224 267028
rect 385276 267016 385282 267028
rect 488534 267016 488540 267028
rect 385276 266988 488540 267016
rect 385276 266976 385282 266988
rect 488534 266976 488540 266988
rect 488592 266976 488598 267028
rect 168466 265616 168472 265668
rect 168524 265656 168530 265668
rect 287238 265656 287244 265668
rect 168524 265628 287244 265656
rect 168524 265616 168530 265628
rect 287238 265616 287244 265628
rect 287296 265616 287302 265668
rect 386414 265616 386420 265668
rect 386472 265656 386478 265668
rect 491294 265656 491300 265668
rect 386472 265628 491300 265656
rect 386472 265616 386478 265628
rect 491294 265616 491300 265628
rect 491352 265616 491358 265668
rect 172514 264188 172520 264240
rect 172572 264228 172578 264240
rect 287146 264228 287152 264240
rect 172572 264200 287152 264228
rect 172572 264188 172578 264200
rect 287146 264188 287152 264200
rect 287204 264188 287210 264240
rect 387978 264188 387984 264240
rect 388036 264228 388042 264240
rect 495434 264228 495440 264240
rect 388036 264200 495440 264228
rect 388036 264188 388042 264200
rect 495434 264188 495440 264200
rect 495492 264188 495498 264240
rect 183554 262828 183560 262880
rect 183612 262868 183618 262880
rect 291286 262868 291292 262880
rect 183612 262840 291292 262868
rect 183612 262828 183618 262840
rect 291286 262828 291292 262840
rect 291344 262828 291350 262880
rect 389174 262828 389180 262880
rect 389232 262868 389238 262880
rect 498286 262868 498292 262880
rect 389232 262840 498292 262868
rect 389232 262828 389238 262840
rect 498286 262828 498292 262840
rect 498344 262828 498350 262880
rect 292574 261536 292580 261588
rect 292632 261576 292638 261588
rect 324590 261576 324596 261588
rect 292632 261548 324596 261576
rect 292632 261536 292638 261548
rect 324590 261536 324596 261548
rect 324648 261536 324654 261588
rect 186314 261468 186320 261520
rect 186372 261508 186378 261520
rect 292758 261508 292764 261520
rect 186372 261480 292764 261508
rect 186372 261468 186378 261480
rect 292758 261468 292764 261480
rect 292816 261468 292822 261520
rect 354858 261468 354864 261520
rect 354916 261508 354922 261520
rect 389174 261508 389180 261520
rect 354916 261480 389180 261508
rect 354916 261468 354922 261480
rect 389174 261468 389180 261480
rect 389232 261468 389238 261520
rect 389358 261468 389364 261520
rect 389416 261508 389422 261520
rect 502334 261508 502340 261520
rect 389416 261480 502340 261508
rect 389416 261468 389422 261480
rect 502334 261468 502340 261480
rect 502392 261468 502398 261520
rect 190454 260108 190460 260160
rect 190512 260148 190518 260160
rect 292850 260148 292856 260160
rect 190512 260120 292856 260148
rect 190512 260108 190518 260120
rect 292850 260108 292856 260120
rect 292908 260108 292914 260160
rect 356238 260108 356244 260160
rect 356296 260148 356302 260160
rect 391934 260148 391940 260160
rect 356296 260120 391940 260148
rect 356296 260108 356302 260120
rect 391934 260108 391940 260120
rect 391992 260108 391998 260160
rect 392118 260108 392124 260160
rect 392176 260148 392182 260160
rect 509234 260148 509240 260160
rect 392176 260120 509240 260148
rect 392176 260108 392182 260120
rect 509234 260108 509240 260120
rect 509292 260108 509298 260160
rect 443638 259360 443644 259412
rect 443696 259400 443702 259412
rect 580166 259400 580172 259412
rect 443696 259372 580172 259400
rect 443696 259360 443702 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 193306 258748 193312 258800
rect 193364 258788 193370 258800
rect 294138 258788 294144 258800
rect 193364 258760 294144 258788
rect 193364 258748 193370 258760
rect 294138 258748 294144 258760
rect 294196 258748 294202 258800
rect 24118 258680 24124 258732
rect 24176 258720 24182 258732
rect 238938 258720 238944 258732
rect 24176 258692 238944 258720
rect 24176 258680 24182 258692
rect 238938 258680 238944 258692
rect 238996 258680 239002 258732
rect 364518 258680 364524 258732
rect 364576 258720 364582 258732
rect 420914 258720 420920 258732
rect 364576 258692 420920 258720
rect 364576 258680 364582 258692
rect 420914 258680 420920 258692
rect 420972 258680 420978 258732
rect 204254 257388 204260 257440
rect 204312 257428 204318 257440
rect 298186 257428 298192 257440
rect 204312 257400 298192 257428
rect 204312 257388 204318 257400
rect 298186 257388 298192 257400
rect 298244 257388 298250 257440
rect 22094 257320 22100 257372
rect 22152 257360 22158 257372
rect 241698 257360 241704 257372
rect 22152 257332 241704 257360
rect 22152 257320 22158 257332
rect 241698 257320 241704 257332
rect 241756 257320 241762 257372
rect 393406 257320 393412 257372
rect 393464 257360 393470 257372
rect 516134 257360 516140 257372
rect 393464 257332 516140 257360
rect 393464 257320 393470 257332
rect 516134 257320 516140 257332
rect 516192 257320 516198 257372
rect 208394 256028 208400 256080
rect 208452 256068 208458 256080
rect 298370 256068 298376 256080
rect 208452 256040 298376 256068
rect 208452 256028 208458 256040
rect 298370 256028 298376 256040
rect 298428 256028 298434 256080
rect 17954 255960 17960 256012
rect 18012 256000 18018 256012
rect 240318 256000 240324 256012
rect 18012 255972 240324 256000
rect 18012 255960 18018 255972
rect 240318 255960 240324 255972
rect 240376 255960 240382 256012
rect 357618 255960 357624 256012
rect 357676 256000 357682 256012
rect 397454 256000 397460 256012
rect 357676 255972 397460 256000
rect 357676 255960 357682 255972
rect 397454 255960 397460 255972
rect 397512 255960 397518 256012
rect 400858 255960 400864 256012
rect 400916 256000 400922 256012
rect 531314 256000 531320 256012
rect 400916 255972 531320 256000
rect 400916 255960 400922 255972
rect 531314 255960 531320 255972
rect 531372 255960 531378 256012
rect 3326 255212 3332 255264
rect 3384 255252 3390 255264
rect 31018 255252 31024 255264
rect 3384 255224 31024 255252
rect 3384 255212 3390 255224
rect 31018 255212 31024 255224
rect 31076 255212 31082 255264
rect 299474 254736 299480 254788
rect 299532 254776 299538 254788
rect 327350 254776 327356 254788
rect 299532 254748 327356 254776
rect 299532 254736 299538 254748
rect 327350 254736 327356 254748
rect 327408 254736 327414 254788
rect 211154 254600 211160 254652
rect 211212 254640 211218 254652
rect 299750 254640 299756 254652
rect 211212 254612 299756 254640
rect 211212 254600 211218 254612
rect 299750 254600 299756 254612
rect 299808 254600 299814 254652
rect 34514 254532 34520 254584
rect 34572 254572 34578 254584
rect 245838 254572 245844 254584
rect 34572 254544 245844 254572
rect 34572 254532 34578 254544
rect 245838 254532 245844 254544
rect 245896 254532 245902 254584
rect 357526 254532 357532 254584
rect 357584 254572 357590 254584
rect 398926 254572 398932 254584
rect 357584 254544 398932 254572
rect 357584 254532 357590 254544
rect 398926 254532 398932 254544
rect 398984 254532 398990 254584
rect 399018 254532 399024 254584
rect 399076 254572 399082 254584
rect 534074 254572 534080 254584
rect 399076 254544 534080 254572
rect 399076 254532 399082 254544
rect 534074 254532 534080 254544
rect 534132 254532 534138 254584
rect 303614 253376 303620 253428
rect 303672 253416 303678 253428
rect 328730 253416 328736 253428
rect 303672 253388 328736 253416
rect 303672 253376 303678 253388
rect 328730 253376 328736 253388
rect 328788 253376 328794 253428
rect 226426 253240 226432 253292
rect 226484 253280 226490 253292
rect 303890 253280 303896 253292
rect 226484 253252 303896 253280
rect 226484 253240 226490 253252
rect 303890 253240 303896 253252
rect 303948 253240 303954 253292
rect 33134 253172 33140 253224
rect 33192 253212 33198 253224
rect 244458 253212 244464 253224
rect 33192 253184 244464 253212
rect 33192 253172 33198 253184
rect 244458 253172 244464 253184
rect 244516 253172 244522 253224
rect 358998 253172 359004 253224
rect 359056 253212 359062 253224
rect 400306 253212 400312 253224
rect 359056 253184 400312 253212
rect 359056 253172 359062 253184
rect 400306 253172 400312 253184
rect 400364 253172 400370 253224
rect 400398 253172 400404 253224
rect 400456 253212 400462 253224
rect 538214 253212 538220 253224
rect 400456 253184 538220 253212
rect 400456 253172 400462 253184
rect 538214 253172 538220 253184
rect 538272 253172 538278 253224
rect 229094 251880 229100 251932
rect 229152 251920 229158 251932
rect 305086 251920 305092 251932
rect 229152 251892 305092 251920
rect 229152 251880 229158 251892
rect 305086 251880 305092 251892
rect 305144 251880 305150 251932
rect 28994 251812 29000 251864
rect 29052 251852 29058 251864
rect 243078 251852 243084 251864
rect 29052 251824 243084 251852
rect 29052 251812 29058 251824
rect 243078 251812 243084 251824
rect 243136 251812 243142 251864
rect 403158 251812 403164 251864
rect 403216 251852 403222 251864
rect 545114 251852 545120 251864
rect 403216 251824 545120 251852
rect 403216 251812 403222 251824
rect 545114 251812 545120 251824
rect 545172 251812 545178 251864
rect 276198 250588 276204 250640
rect 276256 250628 276262 250640
rect 318978 250628 318984 250640
rect 276256 250600 318984 250628
rect 276256 250588 276262 250600
rect 318978 250588 318984 250600
rect 319036 250588 319042 250640
rect 133874 250452 133880 250504
rect 133932 250492 133938 250504
rect 276106 250492 276112 250504
rect 133932 250464 276112 250492
rect 133932 250452 133938 250464
rect 276106 250452 276112 250464
rect 276164 250452 276170 250504
rect 404446 250452 404452 250504
rect 404504 250492 404510 250504
rect 547966 250492 547972 250504
rect 404504 250464 547972 250492
rect 404504 250452 404510 250464
rect 547966 250452 547972 250464
rect 548024 250452 548030 250504
rect 233234 249092 233240 249144
rect 233292 249132 233298 249144
rect 306466 249132 306472 249144
rect 233292 249104 306472 249132
rect 233292 249092 233298 249104
rect 306466 249092 306472 249104
rect 306524 249092 306530 249144
rect 16574 249024 16580 249076
rect 16632 249064 16638 249076
rect 233970 249064 233976 249076
rect 16632 249036 233976 249064
rect 16632 249024 16638 249036
rect 233970 249024 233976 249036
rect 234028 249024 234034 249076
rect 409966 249024 409972 249076
rect 410024 249064 410030 249076
rect 569954 249064 569960 249076
rect 410024 249036 569960 249064
rect 410024 249024 410030 249036
rect 569954 249024 569960 249036
rect 570012 249024 570018 249076
rect 140774 247664 140780 247716
rect 140832 247704 140838 247716
rect 277486 247704 277492 247716
rect 140832 247676 277492 247704
rect 140832 247664 140838 247676
rect 277486 247664 277492 247676
rect 277544 247664 277550 247716
rect 367278 247664 367284 247716
rect 367336 247704 367342 247716
rect 432046 247704 432052 247716
rect 367336 247676 432052 247704
rect 367336 247664 367342 247676
rect 432046 247664 432052 247676
rect 432104 247664 432110 247716
rect 143626 246304 143632 246356
rect 143684 246344 143690 246356
rect 278958 246344 278964 246356
rect 143684 246316 278964 246344
rect 143684 246304 143690 246316
rect 278958 246304 278964 246316
rect 279016 246304 279022 246356
rect 385126 246304 385132 246356
rect 385184 246344 385190 246356
rect 485774 246344 485780 246356
rect 385184 246316 485780 246344
rect 385184 246304 385190 246316
rect 485774 246304 485780 246316
rect 485832 246304 485838 246356
rect 422938 245556 422944 245608
rect 422996 245596 423002 245608
rect 580166 245596 580172 245608
rect 422996 245568 580172 245596
rect 422996 245556 423002 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 147674 244876 147680 244928
rect 147732 244916 147738 244928
rect 280246 244916 280252 244928
rect 147732 244888 280252 244916
rect 147732 244876 147738 244888
rect 280246 244876 280252 244888
rect 280304 244876 280310 244928
rect 386506 243584 386512 243636
rect 386564 243624 386570 243636
rect 386564 243596 393314 243624
rect 386564 243584 386570 243596
rect 151814 243516 151820 243568
rect 151872 243556 151878 243568
rect 281626 243556 281632 243568
rect 151872 243528 281632 243556
rect 151872 243516 151878 243528
rect 281626 243516 281632 243528
rect 281684 243516 281690 243568
rect 353478 243516 353484 243568
rect 353536 243556 353542 243568
rect 386414 243556 386420 243568
rect 353536 243528 386420 243556
rect 353536 243516 353542 243528
rect 386414 243516 386420 243528
rect 386472 243516 386478 243568
rect 393286 243556 393314 243596
rect 492674 243556 492680 243568
rect 393286 243528 492680 243556
rect 492674 243516 492680 243528
rect 492732 243516 492738 243568
rect 158714 242156 158720 242208
rect 158772 242196 158778 242208
rect 283006 242196 283012 242208
rect 158772 242168 283012 242196
rect 158772 242156 158778 242168
rect 283006 242156 283012 242168
rect 283064 242156 283070 242208
rect 387886 242156 387892 242208
rect 387944 242196 387950 242208
rect 496814 242196 496820 242208
rect 387944 242168 496820 242196
rect 387944 242156 387950 242168
rect 496814 242156 496820 242168
rect 496872 242156 496878 242208
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 232590 241448 232596 241460
rect 3292 241420 232596 241448
rect 3292 241408 3298 241420
rect 232590 241408 232596 241420
rect 232648 241408 232654 241460
rect 389266 240728 389272 240780
rect 389324 240768 389330 240780
rect 499574 240768 499580 240780
rect 389324 240740 499580 240768
rect 389324 240728 389330 240740
rect 499574 240728 499580 240740
rect 499632 240728 499638 240780
rect 166994 239368 167000 239420
rect 167052 239408 167058 239420
rect 285766 239408 285772 239420
rect 167052 239380 285772 239408
rect 167052 239368 167058 239380
rect 285766 239368 285772 239380
rect 285824 239368 285830 239420
rect 390646 239368 390652 239420
rect 390704 239408 390710 239420
rect 503714 239408 503720 239420
rect 390704 239380 503720 239408
rect 390704 239368 390710 239380
rect 503714 239368 503720 239380
rect 503772 239368 503778 239420
rect 180794 238008 180800 238060
rect 180852 238048 180858 238060
rect 289998 238048 290004 238060
rect 180852 238020 290004 238048
rect 180852 238008 180858 238020
rect 289998 238008 290004 238020
rect 290056 238008 290062 238060
rect 392026 238008 392032 238060
rect 392084 238048 392090 238060
rect 510614 238048 510620 238060
rect 392084 238020 510620 238048
rect 392084 238008 392090 238020
rect 510614 238008 510620 238020
rect 510672 238008 510678 238060
rect 187694 236648 187700 236700
rect 187752 236688 187758 236700
rect 292666 236688 292672 236700
rect 187752 236660 292672 236688
rect 187752 236648 187758 236660
rect 292666 236648 292672 236660
rect 292724 236648 292730 236700
rect 394786 236648 394792 236700
rect 394844 236688 394850 236700
rect 517514 236688 517520 236700
rect 394844 236660 517520 236688
rect 394844 236648 394850 236660
rect 517514 236648 517520 236660
rect 517572 236648 517578 236700
rect 191834 235220 191840 235272
rect 191892 235260 191898 235272
rect 294046 235260 294052 235272
rect 191892 235232 294052 235260
rect 191892 235220 191898 235232
rect 294046 235220 294052 235232
rect 294104 235220 294110 235272
rect 396258 235220 396264 235272
rect 396316 235260 396322 235272
rect 521654 235260 521660 235272
rect 396316 235232 521660 235260
rect 396316 235220 396322 235232
rect 521654 235220 521660 235232
rect 521712 235220 521718 235272
rect 131114 233860 131120 233912
rect 131172 233900 131178 233912
rect 274726 233900 274732 233912
rect 131172 233872 274732 233900
rect 131172 233860 131178 233872
rect 274726 233860 274732 233872
rect 274784 233860 274790 233912
rect 396166 233860 396172 233912
rect 396224 233900 396230 233912
rect 524414 233900 524420 233912
rect 396224 233872 524420 233900
rect 396224 233860 396230 233872
rect 524414 233860 524420 233872
rect 524472 233860 524478 233912
rect 438118 233180 438124 233232
rect 438176 233220 438182 233232
rect 579614 233220 579620 233232
rect 438176 233192 579620 233220
rect 438176 233180 438182 233192
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 201586 232500 201592 232552
rect 201644 232540 201650 232552
rect 296806 232540 296812 232552
rect 201644 232512 296812 232540
rect 201644 232500 201650 232512
rect 296806 232500 296812 232512
rect 296864 232500 296870 232552
rect 209866 231072 209872 231124
rect 209924 231112 209930 231124
rect 299658 231112 299664 231124
rect 209924 231084 299664 231112
rect 209924 231072 209930 231084
rect 299658 231072 299664 231084
rect 299716 231072 299722 231124
rect 401778 231072 401784 231124
rect 401836 231112 401842 231124
rect 539594 231112 539600 231124
rect 401836 231084 539600 231112
rect 401836 231072 401842 231084
rect 539594 231072 539600 231084
rect 539652 231072 539658 231124
rect 212534 229712 212540 229764
rect 212592 229752 212598 229764
rect 299566 229752 299572 229764
rect 212592 229724 299572 229752
rect 212592 229712 212598 229724
rect 299566 229712 299572 229724
rect 299624 229712 299630 229764
rect 401686 229712 401692 229764
rect 401744 229752 401750 229764
rect 542354 229752 542360 229764
rect 401744 229724 542360 229752
rect 401744 229712 401750 229724
rect 542354 229712 542360 229724
rect 542412 229712 542418 229764
rect 142154 228352 142160 228404
rect 142212 228392 142218 228404
rect 278866 228392 278872 228404
rect 142212 228364 278872 228392
rect 142212 228352 142218 228364
rect 278866 228352 278872 228364
rect 278924 228352 278930 228404
rect 403066 228352 403072 228404
rect 403124 228392 403130 228404
rect 546494 228392 546500 228404
rect 403124 228364 546500 228392
rect 403124 228352 403130 228364
rect 546494 228352 546500 228364
rect 546552 228352 546558 228404
rect 100754 226992 100760 227044
rect 100812 227032 100818 227044
rect 265158 227032 265164 227044
rect 100812 227004 265164 227032
rect 100812 226992 100818 227004
rect 265158 226992 265164 227004
rect 265216 226992 265222 227044
rect 405826 226992 405832 227044
rect 405884 227032 405890 227044
rect 553394 227032 553400 227044
rect 405884 227004 553400 227032
rect 405884 226992 405890 227004
rect 553394 226992 553400 227004
rect 553452 226992 553458 227044
rect 103514 225564 103520 225616
rect 103572 225604 103578 225616
rect 266538 225604 266544 225616
rect 103572 225576 266544 225604
rect 103572 225564 103578 225576
rect 266538 225564 266544 225576
rect 266596 225564 266602 225616
rect 407206 225564 407212 225616
rect 407264 225604 407270 225616
rect 560294 225604 560300 225616
rect 407264 225576 560300 225604
rect 407264 225564 407270 225576
rect 560294 225564 560300 225576
rect 560352 225564 560358 225616
rect 44174 224204 44180 224256
rect 44232 224244 44238 224256
rect 248598 224244 248604 224256
rect 44232 224216 248604 224244
rect 44232 224204 44238 224216
rect 248598 224204 248604 224216
rect 248656 224204 248662 224256
rect 411346 224204 411352 224256
rect 411404 224244 411410 224256
rect 574094 224244 574100 224256
rect 411404 224216 574100 224244
rect 411404 224204 411410 224216
rect 574094 224204 574100 224216
rect 574152 224204 574158 224256
rect 13078 222844 13084 222896
rect 13136 222884 13142 222896
rect 237558 222884 237564 222896
rect 13136 222856 237564 222884
rect 13136 222844 13142 222856
rect 237558 222844 237564 222856
rect 237616 222844 237622 222896
rect 48314 221416 48320 221468
rect 48372 221456 48378 221468
rect 249978 221456 249984 221468
rect 48372 221428 249984 221456
rect 48372 221416 48378 221428
rect 249978 221416 249984 221428
rect 250036 221416 250042 221468
rect 52454 220056 52460 220108
rect 52512 220096 52518 220108
rect 249886 220096 249892 220108
rect 52512 220068 249892 220096
rect 52512 220056 52518 220068
rect 249886 220056 249892 220068
rect 249944 220056 249950 220108
rect 442258 219376 442264 219428
rect 442316 219416 442322 219428
rect 580166 219416 580172 219428
rect 442316 219388 580172 219416
rect 442316 219376 442322 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 59354 218696 59360 218748
rect 59412 218736 59418 218748
rect 252738 218736 252744 218748
rect 59412 218708 252744 218736
rect 59412 218696 59418 218708
rect 252738 218696 252744 218708
rect 252796 218696 252802 218748
rect 62114 217268 62120 217320
rect 62172 217308 62178 217320
rect 251818 217308 251824 217320
rect 62172 217280 251824 217308
rect 62172 217268 62178 217280
rect 251818 217268 251824 217280
rect 251876 217268 251882 217320
rect 66254 215908 66260 215960
rect 66312 215948 66318 215960
rect 255498 215948 255504 215960
rect 66312 215920 255504 215948
rect 66312 215908 66318 215920
rect 255498 215908 255504 215920
rect 255556 215908 255562 215960
rect 2774 214956 2780 215008
rect 2832 214996 2838 215008
rect 4890 214996 4896 215008
rect 2832 214968 4896 214996
rect 2832 214956 2838 214968
rect 4890 214956 4896 214968
rect 4948 214956 4954 215008
rect 84194 214548 84200 214600
rect 84252 214588 84258 214600
rect 261018 214588 261024 214600
rect 84252 214560 261024 214588
rect 84252 214548 84258 214560
rect 261018 214548 261024 214560
rect 261076 214548 261082 214600
rect 86954 213188 86960 213240
rect 87012 213228 87018 213240
rect 260926 213228 260932 213240
rect 87012 213200 260932 213228
rect 87012 213188 87018 213200
rect 260926 213188 260932 213200
rect 260984 213188 260990 213240
rect 97994 211760 98000 211812
rect 98052 211800 98058 211812
rect 265066 211800 265072 211812
rect 98052 211772 265072 211800
rect 98052 211760 98058 211772
rect 265066 211760 265072 211772
rect 265124 211760 265130 211812
rect 104894 210400 104900 210452
rect 104952 210440 104958 210452
rect 266446 210440 266452 210452
rect 104952 210412 266452 210440
rect 104952 210400 104958 210412
rect 266446 210400 266452 210412
rect 266504 210400 266510 210452
rect 30374 209040 30380 209092
rect 30432 209080 30438 209092
rect 244366 209080 244372 209092
rect 30432 209052 244372 209080
rect 30432 209040 30438 209052
rect 244366 209040 244372 209052
rect 244424 209040 244430 209092
rect 41414 207612 41420 207664
rect 41472 207652 41478 207664
rect 247218 207652 247224 207664
rect 41472 207624 247224 207652
rect 41472 207612 41478 207624
rect 247218 207612 247224 207624
rect 247276 207612 247282 207664
rect 421558 206932 421564 206984
rect 421616 206972 421622 206984
rect 580166 206972 580172 206984
rect 421616 206944 580172 206972
rect 421616 206932 421622 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 56594 206252 56600 206304
rect 56652 206292 56658 206304
rect 252646 206292 252652 206304
rect 56652 206264 252652 206292
rect 56652 206252 56658 206264
rect 252646 206252 252652 206264
rect 252704 206252 252710 206304
rect 63494 204892 63500 204944
rect 63552 204932 63558 204944
rect 254210 204932 254216 204944
rect 63552 204904 254216 204932
rect 63552 204892 63558 204904
rect 254210 204892 254216 204904
rect 254268 204892 254274 204944
rect 67634 203532 67640 203584
rect 67692 203572 67698 203584
rect 255406 203572 255412 203584
rect 67692 203544 255412 203572
rect 67692 203532 67698 203544
rect 255406 203532 255412 203544
rect 255464 203532 255470 203584
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 11790 202824 11796 202836
rect 3384 202796 11796 202824
rect 3384 202784 3390 202796
rect 11790 202784 11796 202796
rect 11848 202784 11854 202836
rect 70394 202104 70400 202156
rect 70452 202144 70458 202156
rect 256878 202144 256884 202156
rect 70452 202116 256884 202144
rect 70452 202104 70458 202116
rect 256878 202104 256884 202116
rect 256936 202104 256942 202156
rect 77294 200744 77300 200796
rect 77352 200784 77358 200796
rect 258258 200784 258264 200796
rect 77352 200756 258264 200784
rect 77352 200744 77358 200756
rect 258258 200744 258264 200756
rect 258316 200744 258322 200796
rect 88334 199384 88340 199436
rect 88392 199424 88398 199436
rect 262398 199424 262404 199436
rect 88392 199396 262404 199424
rect 88392 199384 88398 199396
rect 262398 199384 262404 199396
rect 262456 199384 262462 199436
rect 92474 197956 92480 198008
rect 92532 197996 92538 198008
rect 262306 197996 262312 198008
rect 92532 197968 262312 197996
rect 92532 197956 92538 197968
rect 262306 197956 262312 197968
rect 262364 197956 262370 198008
rect 95234 196596 95240 196648
rect 95292 196636 95298 196648
rect 263778 196636 263784 196648
rect 95292 196608 263784 196636
rect 95292 196596 95298 196608
rect 263778 196596 263784 196608
rect 263836 196596 263842 196648
rect 106274 195236 106280 195288
rect 106332 195276 106338 195288
rect 267918 195276 267924 195288
rect 106332 195248 267924 195276
rect 106332 195236 106338 195248
rect 267918 195236 267924 195248
rect 267976 195236 267982 195288
rect 429838 193128 429844 193180
rect 429896 193168 429902 193180
rect 580166 193168 580172 193180
rect 429896 193140 580172 193168
rect 429896 193128 429902 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 40678 189020 40684 189032
rect 3200 188992 40684 189020
rect 3200 188980 3206 188992
rect 40678 188980 40684 188992
rect 40736 188980 40742 189032
rect 440878 179324 440884 179376
rect 440936 179364 440942 179376
rect 580166 179364 580172 179376
rect 440936 179336 580172 179364
rect 440936 179324 440942 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 420178 166948 420184 167000
rect 420236 166988 420242 167000
rect 580166 166988 580172 167000
rect 420236 166960 580172 166988
rect 420236 166948 420242 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 229738 164200 229744 164212
rect 3384 164172 229744 164200
rect 3384 164160 3390 164172
rect 229738 164160 229744 164172
rect 229796 164160 229802 164212
rect 428458 153144 428464 153196
rect 428516 153184 428522 153196
rect 580166 153184 580172 153196
rect 428516 153156 580172 153184
rect 428516 153144 428522 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 13170 150396 13176 150408
rect 3384 150368 13176 150396
rect 3384 150356 3390 150368
rect 13170 150356 13176 150368
rect 13228 150356 13234 150408
rect 439498 139340 439504 139392
rect 439556 139380 439562 139392
rect 580166 139380 580172 139392
rect 439556 139352 580172 139380
rect 439556 139340 439562 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 435358 126896 435364 126948
rect 435416 126936 435422 126948
rect 579614 126936 579620 126948
rect 435416 126908 579620 126936
rect 435416 126896 435422 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 427078 113092 427084 113144
rect 427136 113132 427142 113144
rect 580166 113132 580172 113144
rect 427136 113104 580172 113132
rect 427136 113092 427142 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 7650 111052 7656 111104
rect 7708 111092 7714 111104
rect 234798 111092 234804 111104
rect 7708 111064 234804 111092
rect 7708 111052 7714 111064
rect 234798 111052 234804 111064
rect 234856 111052 234862 111104
rect 3234 110984 3240 111036
rect 3292 111024 3298 111036
rect 7558 111024 7564 111036
rect 3292 110996 7564 111024
rect 3292 110984 3298 110996
rect 7558 110984 7564 110996
rect 7616 110984 7622 111036
rect 436738 100648 436744 100700
rect 436796 100688 436802 100700
rect 579706 100688 579712 100700
rect 436796 100660 579712 100688
rect 436796 100648 436802 100660
rect 579706 100648 579712 100660
rect 579764 100648 579770 100700
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 14458 97968 14464 97980
rect 3292 97940 14464 97968
rect 3292 97928 3298 97940
rect 14458 97928 14464 97940
rect 14516 97928 14522 97980
rect 14550 97248 14556 97300
rect 14608 97288 14614 97300
rect 237466 97288 237472 97300
rect 14608 97260 237472 97288
rect 14608 97248 14614 97260
rect 237466 97248 237472 97260
rect 237524 97248 237530 97300
rect 418798 86912 418804 86964
rect 418856 86952 418862 86964
rect 579982 86952 579988 86964
rect 418856 86924 579988 86952
rect 418856 86912 418862 86924
rect 579982 86912 579988 86924
rect 580040 86912 580046 86964
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 21358 85524 21364 85536
rect 3384 85496 21364 85524
rect 3384 85484 3390 85496
rect 21358 85484 21364 85496
rect 21416 85484 21422 85536
rect 425698 73108 425704 73160
rect 425756 73148 425762 73160
rect 580166 73148 580172 73160
rect 425756 73120 580172 73148
rect 425756 73108 425762 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 233878 71720 233884 71732
rect 3384 71692 233884 71720
rect 3384 71680 3390 71692
rect 233878 71680 233884 71692
rect 233936 71680 233942 71732
rect 27614 68280 27620 68332
rect 27672 68320 27678 68332
rect 242986 68320 242992 68332
rect 27672 68292 242992 68320
rect 27672 68280 27678 68292
rect 242986 68280 242992 68292
rect 243044 68280 243050 68332
rect 44266 64132 44272 64184
rect 44324 64172 44330 64184
rect 248506 64172 248512 64184
rect 44324 64144 248512 64172
rect 44324 64132 44330 64144
rect 248506 64132 248512 64144
rect 248564 64132 248570 64184
rect 99374 62772 99380 62824
rect 99432 62812 99438 62824
rect 265250 62812 265256 62824
rect 99432 62784 265256 62812
rect 99432 62772 99438 62784
rect 265250 62772 265256 62784
rect 265308 62772 265314 62824
rect 52546 61344 52552 61396
rect 52604 61384 52610 61396
rect 251266 61384 251272 61396
rect 52604 61356 251272 61384
rect 52604 61344 52610 61356
rect 251266 61344 251272 61356
rect 251324 61344 251330 61396
rect 432598 60664 432604 60716
rect 432656 60704 432662 60716
rect 579798 60704 579804 60716
rect 432656 60676 579804 60704
rect 432656 60664 432662 60676
rect 579798 60664 579804 60676
rect 579856 60664 579862 60716
rect 102226 59984 102232 60036
rect 102284 60024 102290 60036
rect 266630 60024 266636 60036
rect 102284 59996 266636 60024
rect 102284 59984 102290 59996
rect 266630 59984 266636 59996
rect 266688 59984 266694 60036
rect 3326 59304 3332 59356
rect 3384 59344 3390 59356
rect 28258 59344 28264 59356
rect 3384 59316 28264 59344
rect 3384 59304 3390 59316
rect 28258 59304 28264 59316
rect 28316 59304 28322 59356
rect 160186 58624 160192 58676
rect 160244 58664 160250 58676
rect 284386 58664 284392 58676
rect 160244 58636 284392 58664
rect 160244 58624 160250 58636
rect 284386 58624 284392 58636
rect 284444 58624 284450 58676
rect 155954 57196 155960 57248
rect 156012 57236 156018 57248
rect 282914 57236 282920 57248
rect 156012 57208 282920 57236
rect 156012 57196 156018 57208
rect 282914 57196 282920 57208
rect 282972 57196 282978 57248
rect 151906 55836 151912 55888
rect 151964 55876 151970 55888
rect 281534 55876 281540 55888
rect 151964 55848 281540 55876
rect 151964 55836 151970 55848
rect 281534 55836 281540 55848
rect 281592 55836 281598 55888
rect 135346 54476 135352 54528
rect 135404 54516 135410 54528
rect 276014 54516 276020 54528
rect 135404 54488 276020 54516
rect 135404 54476 135410 54488
rect 276014 54476 276020 54488
rect 276072 54476 276078 54528
rect 149054 53048 149060 53100
rect 149112 53088 149118 53100
rect 280154 53088 280160 53100
rect 149112 53060 280160 53088
rect 149112 53048 149118 53060
rect 280154 53048 280160 53060
rect 280212 53048 280218 53100
rect 69106 51688 69112 51740
rect 69164 51728 69170 51740
rect 255314 51728 255320 51740
rect 69164 51700 255320 51728
rect 69164 51688 69170 51700
rect 255314 51688 255320 51700
rect 255372 51688 255378 51740
rect 255406 51688 255412 51740
rect 255464 51728 255470 51740
rect 313366 51728 313372 51740
rect 255464 51700 313372 51728
rect 255464 51688 255470 51700
rect 313366 51688 313372 51700
rect 313424 51688 313430 51740
rect 396074 51688 396080 51740
rect 396132 51728 396138 51740
rect 523034 51728 523040 51740
rect 396132 51700 523040 51728
rect 396132 51688 396138 51700
rect 523034 51688 523040 51700
rect 523092 51688 523098 51740
rect 49694 50328 49700 50380
rect 49752 50368 49758 50380
rect 249794 50368 249800 50380
rect 49752 50340 249800 50368
rect 49752 50328 49758 50340
rect 249794 50328 249800 50340
rect 249852 50328 249858 50380
rect 251266 50328 251272 50380
rect 251324 50368 251330 50380
rect 312078 50368 312084 50380
rect 251324 50340 312084 50368
rect 251324 50328 251330 50340
rect 312078 50328 312084 50340
rect 312136 50328 312142 50380
rect 244366 48968 244372 49020
rect 244424 49008 244430 49020
rect 310698 49008 310704 49020
rect 244424 48980 310704 49008
rect 244424 48968 244430 48980
rect 310698 48968 310704 48980
rect 310756 48968 310762 49020
rect 237466 47540 237472 47592
rect 237524 47580 237530 47592
rect 307846 47580 307852 47592
rect 237524 47552 307852 47580
rect 237524 47540 237530 47552
rect 307846 47540 307852 47552
rect 307904 47540 307910 47592
rect 417418 46860 417424 46912
rect 417476 46900 417482 46912
rect 580166 46900 580172 46912
rect 417476 46872 580172 46900
rect 417476 46860 417482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 234614 46180 234620 46232
rect 234672 46220 234678 46232
rect 305638 46220 305644 46232
rect 234672 46192 305644 46220
rect 234672 46180 234678 46192
rect 305638 46180 305644 46192
rect 305696 46180 305702 46232
rect 363138 46180 363144 46232
rect 363196 46220 363202 46232
rect 416774 46220 416780 46232
rect 363196 46192 416780 46220
rect 363196 46180 363202 46192
rect 416774 46180 416780 46192
rect 416832 46180 416838 46232
rect 230474 44820 230480 44872
rect 230532 44860 230538 44872
rect 304994 44860 305000 44872
rect 230532 44832 305000 44860
rect 230532 44820 230538 44832
rect 304994 44820 305000 44832
rect 305052 44820 305058 44872
rect 216674 43392 216680 43444
rect 216732 43432 216738 43444
rect 300854 43432 300860 43444
rect 216732 43404 300860 43432
rect 216732 43392 216738 43404
rect 300854 43392 300860 43404
rect 300912 43392 300918 43444
rect 198734 42032 198740 42084
rect 198792 42072 198798 42084
rect 295426 42072 295432 42084
rect 198792 42044 295432 42072
rect 198792 42032 198798 42044
rect 295426 42032 295432 42044
rect 295484 42032 295490 42084
rect 194594 40672 194600 40724
rect 194652 40712 194658 40724
rect 294230 40712 294236 40724
rect 194652 40684 294236 40712
rect 194652 40672 194658 40684
rect 294230 40672 294236 40684
rect 294288 40672 294294 40724
rect 185026 39312 185032 39364
rect 185084 39352 185090 39364
rect 291470 39352 291476 39364
rect 185084 39324 291476 39352
rect 185084 39312 185090 39324
rect 291470 39312 291476 39324
rect 291528 39312 291534 39364
rect 310698 39312 310704 39364
rect 310756 39352 310762 39364
rect 330110 39352 330116 39364
rect 310756 39324 330116 39352
rect 310756 39312 310762 39324
rect 330110 39312 330116 39324
rect 330168 39312 330174 39364
rect 169754 37884 169760 37936
rect 169812 37924 169818 37936
rect 287330 37924 287336 37936
rect 169812 37896 287336 37924
rect 169812 37884 169818 37896
rect 287330 37884 287336 37896
rect 287388 37884 287394 37936
rect 138014 36524 138020 36576
rect 138072 36564 138078 36576
rect 277670 36564 277676 36576
rect 138072 36536 277676 36564
rect 138072 36524 138078 36536
rect 277670 36524 277676 36536
rect 277728 36524 277734 36576
rect 282914 36524 282920 36576
rect 282972 36564 282978 36576
rect 321830 36564 321836 36576
rect 282972 36536 321836 36564
rect 282972 36524 282978 36536
rect 321830 36524 321836 36536
rect 321888 36524 321894 36576
rect 85666 35164 85672 35216
rect 85724 35204 85730 35216
rect 260834 35204 260840 35216
rect 85724 35176 260840 35204
rect 85724 35164 85730 35176
rect 260834 35164 260840 35176
rect 260892 35164 260898 35216
rect 267918 35164 267924 35216
rect 267976 35204 267982 35216
rect 317598 35204 317604 35216
rect 267976 35176 317604 35204
rect 267976 35164 267982 35176
rect 317598 35164 317604 35176
rect 317656 35164 317662 35216
rect 73154 33736 73160 33788
rect 73212 33776 73218 33788
rect 256786 33776 256792 33788
rect 73212 33748 256792 33776
rect 73212 33736 73218 33748
rect 256786 33736 256792 33748
rect 256844 33736 256850 33788
rect 258258 33736 258264 33788
rect 258316 33776 258322 33788
rect 314746 33776 314752 33788
rect 258316 33748 314752 33776
rect 258316 33736 258322 33748
rect 314746 33736 314752 33748
rect 314804 33736 314810 33788
rect 2774 32444 2780 32496
rect 2832 32484 2838 32496
rect 6178 32484 6184 32496
rect 2832 32456 6184 32484
rect 2832 32444 2838 32456
rect 6178 32444 6184 32456
rect 6236 32444 6242 32496
rect 55214 32376 55220 32428
rect 55272 32416 55278 32428
rect 251174 32416 251180 32428
rect 55272 32388 251180 32416
rect 55272 32376 55278 32388
rect 251174 32376 251180 32388
rect 251232 32376 251238 32428
rect 251358 32376 251364 32428
rect 251416 32416 251422 32428
rect 311986 32416 311992 32428
rect 251416 32388 311992 32416
rect 251416 32376 251422 32388
rect 311986 32376 311992 32388
rect 312044 32376 312050 32428
rect 358906 32376 358912 32428
rect 358964 32416 358970 32428
rect 404446 32416 404452 32428
rect 358964 32388 404452 32416
rect 358964 32376 358970 32388
rect 404446 32376 404452 32388
rect 404504 32376 404510 32428
rect 411254 32376 411260 32428
rect 411312 32416 411318 32428
rect 571334 32416 571340 32428
rect 411312 32388 571340 32416
rect 411312 32376 411318 32388
rect 571334 32376 571340 32388
rect 571392 32376 571398 32428
rect 247218 31016 247224 31068
rect 247276 31056 247282 31068
rect 310606 31056 310612 31068
rect 247276 31028 310612 31056
rect 247276 31016 247282 31028
rect 310606 31016 310612 31028
rect 310664 31016 310670 31068
rect 356146 31016 356152 31068
rect 356204 31056 356210 31068
rect 393406 31056 393412 31068
rect 356204 31028 393412 31056
rect 356204 31016 356210 31028
rect 393406 31016 393412 31028
rect 393464 31016 393470 31068
rect 242986 29588 242992 29640
rect 243044 29628 243050 29640
rect 309318 29628 309324 29640
rect 243044 29600 309324 29628
rect 243044 29588 243050 29600
rect 309318 29588 309324 29600
rect 309376 29588 309382 29640
rect 354766 29588 354772 29640
rect 354824 29628 354830 29640
rect 390738 29628 390744 29640
rect 354824 29600 390744 29628
rect 354824 29588 354830 29600
rect 390738 29588 390744 29600
rect 390796 29588 390802 29640
rect 400214 29588 400220 29640
rect 400272 29628 400278 29640
rect 535454 29628 535460 29640
rect 400272 29600 535460 29628
rect 400272 29588 400278 29600
rect 535454 29588 535460 29600
rect 535512 29588 535518 29640
rect 240318 28228 240324 28280
rect 240376 28268 240382 28280
rect 309226 28268 309232 28280
rect 240376 28240 309232 28268
rect 240376 28228 240382 28240
rect 309226 28228 309232 28240
rect 309284 28228 309290 28280
rect 350626 28228 350632 28280
rect 350684 28268 350690 28280
rect 375558 28268 375564 28280
rect 350684 28240 375564 28268
rect 350684 28228 350690 28240
rect 375558 28228 375564 28240
rect 375616 28228 375622 28280
rect 393314 28228 393320 28280
rect 393372 28268 393378 28280
rect 514846 28268 514852 28280
rect 393372 28240 514852 28268
rect 393372 28228 393378 28240
rect 514846 28228 514852 28240
rect 514904 28228 514910 28280
rect 262306 26936 262312 26988
rect 262364 26976 262370 26988
rect 316218 26976 316224 26988
rect 262364 26948 316224 26976
rect 262364 26936 262370 26948
rect 316218 26936 316224 26948
rect 316276 26936 316282 26988
rect 218054 26868 218060 26920
rect 218112 26908 218118 26920
rect 298738 26908 298744 26920
rect 218112 26880 298744 26908
rect 218112 26868 218118 26880
rect 298738 26868 298744 26880
rect 298796 26868 298802 26920
rect 347958 26868 347964 26920
rect 348016 26908 348022 26920
rect 365806 26908 365812 26920
rect 348016 26880 365812 26908
rect 348016 26868 348022 26880
rect 365806 26868 365812 26880
rect 365864 26868 365870 26920
rect 390554 26868 390560 26920
rect 390612 26908 390618 26920
rect 506566 26908 506572 26920
rect 390612 26880 506572 26908
rect 390612 26868 390618 26880
rect 506566 26868 506572 26880
rect 506624 26868 506630 26920
rect 162854 25576 162860 25628
rect 162912 25616 162918 25628
rect 284570 25616 284576 25628
rect 162912 25588 284576 25616
rect 162912 25576 162918 25588
rect 284570 25576 284576 25588
rect 284628 25576 284634 25628
rect 284386 25508 284392 25560
rect 284444 25548 284450 25560
rect 323118 25548 323124 25560
rect 284444 25520 323124 25548
rect 284444 25508 284450 25520
rect 323118 25508 323124 25520
rect 323176 25508 323182 25560
rect 360378 25508 360384 25560
rect 360436 25548 360442 25560
rect 407206 25548 407212 25560
rect 360436 25520 407212 25548
rect 360436 25508 360442 25520
rect 407206 25508 407212 25520
rect 407264 25508 407270 25560
rect 408494 25508 408500 25560
rect 408552 25548 408558 25560
rect 564526 25548 564532 25560
rect 408552 25520 564532 25548
rect 408552 25508 408558 25520
rect 564526 25508 564532 25520
rect 564584 25508 564590 25560
rect 353386 24216 353392 24268
rect 353444 24256 353450 24268
rect 385126 24256 385132 24268
rect 353444 24228 385132 24256
rect 353444 24216 353450 24228
rect 385126 24216 385132 24228
rect 385184 24216 385190 24268
rect 259730 24148 259736 24200
rect 259788 24188 259794 24200
rect 307110 24188 307116 24200
rect 259788 24160 307116 24188
rect 259788 24148 259794 24160
rect 307110 24148 307116 24160
rect 307168 24148 307174 24200
rect 126974 24080 126980 24132
rect 127032 24120 127038 24132
rect 273346 24120 273352 24132
rect 127032 24092 273352 24120
rect 127032 24080 127038 24092
rect 273346 24080 273352 24092
rect 273404 24080 273410 24132
rect 281534 24080 281540 24132
rect 281592 24120 281598 24132
rect 321738 24120 321744 24132
rect 281592 24092 321744 24120
rect 281592 24080 281598 24092
rect 321738 24080 321744 24092
rect 321796 24080 321802 24132
rect 385034 24080 385040 24132
rect 385092 24120 385098 24132
rect 490006 24120 490012 24132
rect 385092 24092 490012 24120
rect 385092 24080 385098 24092
rect 490006 24080 490012 24092
rect 490064 24080 490070 24132
rect 248506 22788 248512 22840
rect 248564 22828 248570 22840
rect 310790 22828 310796 22840
rect 248564 22800 310796 22828
rect 248564 22788 248570 22800
rect 310790 22788 310796 22800
rect 310848 22788 310854 22840
rect 60826 22720 60832 22772
rect 60884 22760 60890 22772
rect 252830 22760 252836 22772
rect 60884 22732 252836 22760
rect 60884 22720 60890 22732
rect 252830 22720 252836 22732
rect 252888 22720 252894 22772
rect 263778 22720 263784 22772
rect 263836 22760 263842 22772
rect 316126 22760 316132 22772
rect 263836 22732 316132 22760
rect 263836 22720 263842 22732
rect 316126 22720 316132 22732
rect 316184 22720 316190 22772
rect 356054 22720 356060 22772
rect 356112 22760 356118 22772
rect 396074 22760 396080 22772
rect 356112 22732 396080 22760
rect 356112 22720 356118 22732
rect 396074 22720 396080 22732
rect 396132 22720 396138 22772
rect 398834 22720 398840 22772
rect 398892 22760 398898 22772
rect 531406 22760 531412 22772
rect 398892 22732 531412 22760
rect 398892 22720 398898 22732
rect 531406 22720 531412 22732
rect 531464 22720 531470 22772
rect 256786 21428 256792 21480
rect 256844 21468 256850 21480
rect 313458 21468 313464 21480
rect 256844 21440 313464 21468
rect 256844 21428 256850 21440
rect 313458 21428 313464 21440
rect 313516 21428 313522 21480
rect 144914 21360 144920 21412
rect 144972 21400 144978 21412
rect 278774 21400 278780 21412
rect 144972 21372 278780 21400
rect 144972 21360 144978 21372
rect 278774 21360 278780 21372
rect 278832 21360 278838 21412
rect 352098 21360 352104 21412
rect 352156 21400 352162 21412
rect 382458 21400 382464 21412
rect 352156 21372 382464 21400
rect 352156 21360 352162 21372
rect 382458 21360 382464 21372
rect 382516 21360 382522 21412
rect 383654 21360 383660 21412
rect 383712 21400 383718 21412
rect 481726 21400 481732 21412
rect 383712 21372 481732 21400
rect 383712 21360 383718 21372
rect 481726 21360 481732 21372
rect 481784 21360 481790 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 414934 20652 414940 20664
rect 3568 20624 414940 20652
rect 3568 20612 3574 20624
rect 414934 20612 414940 20624
rect 414992 20612 414998 20664
rect 360286 18708 360292 18760
rect 360344 18748 360350 18760
rect 405826 18748 405832 18760
rect 360344 18720 405832 18748
rect 360344 18708 360350 18720
rect 405826 18708 405832 18720
rect 405884 18708 405890 18760
rect 289814 18640 289820 18692
rect 289872 18680 289878 18692
rect 315298 18680 315304 18692
rect 289872 18652 315304 18680
rect 289872 18640 289878 18652
rect 315298 18640 315304 18652
rect 315356 18640 315362 18692
rect 37274 18572 37280 18624
rect 37332 18612 37338 18624
rect 245746 18612 245752 18624
rect 37332 18584 245752 18612
rect 37332 18572 37338 18584
rect 245746 18572 245752 18584
rect 245804 18572 245810 18624
rect 249794 18572 249800 18624
rect 249852 18612 249858 18624
rect 297358 18612 297364 18624
rect 249852 18584 297364 18612
rect 249852 18572 249858 18584
rect 297358 18572 297364 18584
rect 297416 18572 297422 18624
rect 405734 18572 405740 18624
rect 405792 18612 405798 18624
rect 556246 18612 556252 18624
rect 405792 18584 556252 18612
rect 405792 18572 405798 18584
rect 556246 18572 556252 18584
rect 556304 18572 556310 18624
rect 243078 17280 243084 17332
rect 243136 17320 243142 17332
rect 302970 17320 302976 17332
rect 243136 17292 302976 17320
rect 243136 17280 243142 17292
rect 302970 17280 302976 17292
rect 303028 17280 303034 17332
rect 358078 17280 358084 17332
rect 358136 17320 358142 17332
rect 372798 17320 372804 17332
rect 358136 17292 372804 17320
rect 358136 17280 358142 17292
rect 372798 17280 372804 17292
rect 372856 17280 372862 17332
rect 241698 17212 241704 17264
rect 241756 17252 241762 17264
rect 309410 17252 309416 17264
rect 241756 17224 309416 17252
rect 241756 17212 241762 17224
rect 309410 17212 309416 17224
rect 309468 17212 309474 17264
rect 346578 17212 346584 17264
rect 346636 17252 346642 17264
rect 360286 17252 360292 17264
rect 346636 17224 360292 17252
rect 346636 17212 346642 17224
rect 360286 17212 360292 17224
rect 360344 17212 360350 17264
rect 370498 17212 370504 17264
rect 370556 17252 370562 17264
rect 412818 17252 412824 17264
rect 370556 17224 412824 17252
rect 370556 17212 370562 17224
rect 412818 17212 412824 17224
rect 412876 17212 412882 17264
rect 260650 15920 260656 15972
rect 260708 15960 260714 15972
rect 291838 15960 291844 15972
rect 260708 15932 291844 15960
rect 260708 15920 260714 15932
rect 291838 15920 291844 15932
rect 291896 15920 291902 15972
rect 116394 15852 116400 15904
rect 116452 15892 116458 15904
rect 270678 15892 270684 15904
rect 116452 15864 270684 15892
rect 116452 15852 116458 15864
rect 270678 15852 270684 15864
rect 270736 15852 270742 15904
rect 279050 15852 279056 15904
rect 279108 15892 279114 15904
rect 319438 15892 319444 15904
rect 279108 15864 319444 15892
rect 279108 15852 279114 15864
rect 319438 15852 319444 15864
rect 319496 15852 319502 15904
rect 358814 15852 358820 15904
rect 358872 15892 358878 15904
rect 402514 15892 402520 15904
rect 358872 15864 402520 15892
rect 358872 15852 358878 15864
rect 402514 15852 402520 15864
rect 402572 15852 402578 15904
rect 404354 15852 404360 15904
rect 404412 15892 404418 15904
rect 550266 15892 550272 15904
rect 404412 15864 550272 15892
rect 404412 15852 404418 15864
rect 550266 15852 550272 15864
rect 550324 15852 550330 15904
rect 112346 14764 112352 14816
rect 112404 14804 112410 14816
rect 269298 14804 269304 14816
rect 112404 14776 269304 14804
rect 112404 14764 112410 14776
rect 269298 14764 269304 14776
rect 269356 14764 269362 14816
rect 109034 14696 109040 14748
rect 109092 14736 109098 14748
rect 267826 14736 267832 14748
rect 109092 14708 267832 14736
rect 109092 14696 109098 14708
rect 267826 14696 267832 14708
rect 267884 14696 267890 14748
rect 93854 14628 93860 14680
rect 93912 14668 93918 14680
rect 263686 14668 263692 14680
rect 93912 14640 263692 14668
rect 93912 14628 93918 14640
rect 263686 14628 263692 14640
rect 263744 14628 263750 14680
rect 91554 14560 91560 14612
rect 91612 14600 91618 14612
rect 262214 14600 262220 14612
rect 91612 14572 262220 14600
rect 91612 14560 91618 14572
rect 262214 14560 262220 14572
rect 262272 14560 262278 14612
rect 80882 14492 80888 14544
rect 80940 14532 80946 14544
rect 259638 14532 259644 14544
rect 80940 14504 259644 14532
rect 80940 14492 80946 14504
rect 259638 14492 259644 14504
rect 259696 14492 259702 14544
rect 77386 14424 77392 14476
rect 77444 14464 77450 14476
rect 258166 14464 258172 14476
rect 77444 14436 258172 14464
rect 77444 14424 77450 14436
rect 258166 14424 258172 14436
rect 258224 14424 258230 14476
rect 267734 14424 267740 14476
rect 267792 14464 267798 14476
rect 313918 14464 313924 14476
rect 267792 14436 313924 14464
rect 267792 14424 267798 14436
rect 313918 14424 313924 14436
rect 313976 14424 313982 14476
rect 352006 14424 352012 14476
rect 352064 14464 352070 14476
rect 381170 14464 381176 14476
rect 352064 14436 381176 14464
rect 352064 14424 352070 14436
rect 381170 14424 381176 14436
rect 381228 14424 381234 14476
rect 407114 14424 407120 14476
rect 407172 14464 407178 14476
rect 559282 14464 559288 14476
rect 407172 14436 559288 14464
rect 407172 14424 407178 14436
rect 559282 14424 559288 14436
rect 559340 14424 559346 14476
rect 313826 13948 313832 14000
rect 313884 13988 313890 14000
rect 318058 13988 318064 14000
rect 313884 13960 318064 13988
rect 313884 13948 313890 13960
rect 318058 13948 318064 13960
rect 318116 13948 318122 14000
rect 118786 13336 118792 13388
rect 118844 13376 118850 13388
rect 270586 13376 270592 13388
rect 118844 13348 270592 13376
rect 118844 13336 118850 13348
rect 270586 13336 270592 13348
rect 270644 13336 270650 13388
rect 114738 13268 114744 13320
rect 114796 13308 114802 13320
rect 270770 13308 270776 13320
rect 114796 13280 270776 13308
rect 114796 13268 114802 13280
rect 270770 13268 270776 13280
rect 270828 13268 270834 13320
rect 111610 13200 111616 13252
rect 111668 13240 111674 13252
rect 269206 13240 269212 13252
rect 111668 13212 269212 13240
rect 111668 13200 111674 13212
rect 269206 13200 269212 13212
rect 269264 13200 269270 13252
rect 108114 13132 108120 13184
rect 108172 13172 108178 13184
rect 268102 13172 268108 13184
rect 108172 13144 268108 13172
rect 108172 13132 108178 13144
rect 268102 13132 268108 13144
rect 268160 13132 268166 13184
rect 350534 13132 350540 13184
rect 350592 13172 350598 13184
rect 377306 13172 377312 13184
rect 350592 13144 377312 13172
rect 350592 13132 350598 13144
rect 377306 13132 377312 13144
rect 377364 13132 377370 13184
rect 93946 13064 93952 13116
rect 94004 13104 94010 13116
rect 263594 13104 263600 13116
rect 94004 13076 263600 13104
rect 94004 13064 94010 13076
rect 263594 13064 263600 13076
rect 263652 13064 263658 13116
rect 270770 13064 270776 13116
rect 270828 13104 270834 13116
rect 317506 13104 317512 13116
rect 270828 13076 317512 13104
rect 270828 13064 270834 13076
rect 317506 13064 317512 13076
rect 317564 13064 317570 13116
rect 363046 13064 363052 13116
rect 363104 13104 363110 13116
rect 415486 13104 415492 13116
rect 363104 13076 415492 13104
rect 363104 13064 363110 13076
rect 415486 13064 415492 13076
rect 415544 13064 415550 13116
rect 417510 13064 417516 13116
rect 417568 13104 417574 13116
rect 541986 13104 541992 13116
rect 417568 13076 541992 13104
rect 417568 13064 417574 13076
rect 541986 13064 541992 13076
rect 542044 13064 542050 13116
rect 160094 11772 160100 11824
rect 160152 11812 160158 11824
rect 161290 11812 161296 11824
rect 160152 11784 161296 11812
rect 160152 11772 160158 11784
rect 161290 11772 161296 11784
rect 161348 11772 161354 11824
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 226334 11772 226340 11824
rect 226392 11812 226398 11824
rect 227530 11812 227536 11824
rect 226392 11784 227536 11812
rect 226392 11772 226398 11784
rect 227530 11772 227536 11784
rect 227588 11772 227594 11824
rect 254210 11772 254216 11824
rect 254268 11812 254274 11824
rect 307018 11812 307024 11824
rect 254268 11784 307024 11812
rect 254268 11772 254274 11784
rect 307018 11772 307024 11784
rect 307076 11772 307082 11824
rect 349338 11772 349344 11824
rect 349396 11812 349402 11824
rect 374270 11812 374276 11824
rect 349396 11784 374276 11812
rect 349396 11772 349402 11784
rect 374270 11772 374276 11784
rect 374328 11772 374334 11824
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 238846 11744 238852 11756
rect 13044 11716 238852 11744
rect 13044 11704 13050 11716
rect 238846 11704 238852 11716
rect 238904 11704 238910 11756
rect 239306 11704 239312 11756
rect 239364 11744 239370 11756
rect 301498 11744 301504 11756
rect 239364 11716 301504 11744
rect 239364 11704 239370 11716
rect 301498 11704 301504 11716
rect 301556 11704 301562 11756
rect 307938 11704 307944 11756
rect 307996 11744 308002 11756
rect 330018 11744 330024 11756
rect 307996 11716 330024 11744
rect 307996 11704 308002 11716
rect 330018 11704 330024 11716
rect 330076 11704 330082 11756
rect 373258 11704 373264 11756
rect 373316 11744 373322 11756
rect 414014 11744 414020 11756
rect 373316 11716 414020 11744
rect 373316 11704 373322 11716
rect 414014 11704 414020 11716
rect 414072 11704 414078 11756
rect 424318 11704 424324 11756
rect 424376 11744 424382 11756
rect 523126 11744 523132 11756
rect 424376 11716 523132 11744
rect 424376 11704 424382 11716
rect 523126 11704 523132 11716
rect 523184 11704 523190 11756
rect 372614 10820 372620 10872
rect 372672 10860 372678 10872
rect 445754 10860 445760 10872
rect 372672 10832 445760 10860
rect 372672 10820 372678 10832
rect 445754 10820 445760 10832
rect 445812 10820 445818 10872
rect 372706 10752 372712 10804
rect 372764 10792 372770 10804
rect 448606 10792 448612 10804
rect 372764 10764 448612 10792
rect 372764 10752 372770 10764
rect 448606 10752 448612 10764
rect 448664 10752 448670 10804
rect 374178 10684 374184 10736
rect 374236 10724 374242 10736
rect 453298 10724 453304 10736
rect 374236 10696 453304 10724
rect 374236 10684 374242 10696
rect 453298 10684 453304 10696
rect 453356 10684 453362 10736
rect 375466 10616 375472 10668
rect 375524 10656 375530 10668
rect 456886 10656 456892 10668
rect 375524 10628 456892 10656
rect 375524 10616 375530 10628
rect 456886 10616 456892 10628
rect 456944 10616 456950 10668
rect 376754 10548 376760 10600
rect 376812 10588 376818 10600
rect 459922 10588 459928 10600
rect 376812 10560 459928 10588
rect 376812 10548 376818 10560
rect 459922 10548 459928 10560
rect 459980 10548 459986 10600
rect 378318 10480 378324 10532
rect 378376 10520 378382 10532
rect 463970 10520 463976 10532
rect 378376 10492 463976 10520
rect 378376 10480 378382 10492
rect 463970 10480 463976 10492
rect 464028 10480 464034 10532
rect 173894 10412 173900 10464
rect 173952 10452 173958 10464
rect 288526 10452 288532 10464
rect 173952 10424 288532 10452
rect 173952 10412 173958 10424
rect 288526 10412 288532 10424
rect 288584 10412 288590 10464
rect 378226 10412 378232 10464
rect 378284 10452 378290 10464
rect 467466 10452 467472 10464
rect 378284 10424 467472 10452
rect 378284 10412 378290 10424
rect 467466 10412 467472 10424
rect 467524 10412 467530 10464
rect 83274 10344 83280 10396
rect 83332 10384 83338 10396
rect 259546 10384 259552 10396
rect 83332 10356 259552 10384
rect 83332 10344 83338 10356
rect 259546 10344 259552 10356
rect 259604 10344 259610 10396
rect 288986 10344 288992 10396
rect 289044 10384 289050 10396
rect 323026 10384 323032 10396
rect 289044 10356 323032 10384
rect 289044 10344 289050 10356
rect 323026 10344 323032 10356
rect 323084 10344 323090 10396
rect 345106 10344 345112 10396
rect 345164 10384 345170 10396
rect 357526 10384 357532 10396
rect 345164 10356 357532 10384
rect 345164 10344 345170 10356
rect 357526 10344 357532 10356
rect 357584 10344 357590 10396
rect 380986 10344 380992 10396
rect 381044 10384 381050 10396
rect 474090 10384 474096 10396
rect 381044 10356 474096 10384
rect 381044 10344 381050 10356
rect 474090 10344 474096 10356
rect 474148 10344 474154 10396
rect 79226 10276 79232 10328
rect 79284 10316 79290 10328
rect 259454 10316 259460 10328
rect 79284 10288 259460 10316
rect 79284 10276 79290 10288
rect 259454 10276 259460 10288
rect 259512 10276 259518 10328
rect 264974 10276 264980 10328
rect 265032 10316 265038 10328
rect 302878 10316 302884 10328
rect 265032 10288 302884 10316
rect 265032 10276 265038 10288
rect 302878 10276 302884 10288
rect 302936 10276 302942 10328
rect 349246 10276 349252 10328
rect 349304 10316 349310 10328
rect 371510 10316 371516 10328
rect 349304 10288 371516 10316
rect 349304 10276 349310 10288
rect 371510 10276 371516 10288
rect 371568 10276 371574 10328
rect 382366 10276 382372 10328
rect 382424 10316 382430 10328
rect 478138 10316 478144 10328
rect 382424 10288 478144 10316
rect 382424 10276 382430 10288
rect 478138 10276 478144 10288
rect 478196 10276 478202 10328
rect 209682 9596 209688 9648
rect 209740 9636 209746 9648
rect 210970 9636 210976 9648
rect 209740 9608 210976 9636
rect 209740 9596 209746 9608
rect 210970 9596 210976 9608
rect 211028 9596 211034 9648
rect 253474 9052 253480 9104
rect 253532 9092 253538 9104
rect 312170 9092 312176 9104
rect 253532 9064 312176 9092
rect 253532 9052 253538 9064
rect 312170 9052 312176 9064
rect 312228 9052 312234 9104
rect 76190 8984 76196 9036
rect 76248 9024 76254 9036
rect 258074 9024 258080 9036
rect 76248 8996 258080 9024
rect 76248 8984 76254 8996
rect 258074 8984 258080 8996
rect 258132 8984 258138 9036
rect 349154 8984 349160 9036
rect 349212 9024 349218 9036
rect 370590 9024 370596 9036
rect 349212 8996 370596 9024
rect 349212 8984 349218 8996
rect 370590 8984 370596 8996
rect 370648 8984 370654 9036
rect 72602 8916 72608 8968
rect 72660 8956 72666 8968
rect 256694 8956 256700 8968
rect 72660 8928 256700 8956
rect 72660 8916 72666 8928
rect 256694 8916 256700 8928
rect 256752 8916 256758 8968
rect 261754 8916 261760 8968
rect 261812 8956 261818 8968
rect 314838 8956 314844 8968
rect 261812 8928 314844 8956
rect 261812 8916 261818 8928
rect 314838 8916 314844 8928
rect 314896 8916 314902 8968
rect 317322 8916 317328 8968
rect 317380 8956 317386 8968
rect 332778 8956 332784 8968
rect 317380 8928 332784 8956
rect 317380 8916 317386 8928
rect 332778 8916 332784 8928
rect 332836 8916 332842 8968
rect 351914 8916 351920 8968
rect 351972 8956 351978 8968
rect 379974 8956 379980 8968
rect 351972 8928 379980 8956
rect 351972 8916 351978 8928
rect 379974 8916 379980 8928
rect 380032 8916 380038 8968
rect 387058 8916 387064 8968
rect 387116 8956 387122 8968
rect 398834 8956 398840 8968
rect 387116 8928 398840 8956
rect 387116 8916 387122 8928
rect 398834 8916 398840 8928
rect 398892 8916 398898 8968
rect 412726 8916 412732 8968
rect 412784 8956 412790 8968
rect 577406 8956 577412 8968
rect 412784 8928 577412 8956
rect 412784 8916 412790 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 377398 8236 377404 8288
rect 377456 8276 377462 8288
rect 378870 8276 378876 8288
rect 377456 8248 378876 8276
rect 377456 8236 377462 8248
rect 378870 8236 378876 8248
rect 378928 8236 378934 8288
rect 272426 7692 272432 7744
rect 272484 7732 272490 7744
rect 318886 7732 318892 7744
rect 272484 7704 318892 7732
rect 272484 7692 272490 7704
rect 318886 7692 318892 7704
rect 318944 7692 318950 7744
rect 197906 7624 197912 7676
rect 197964 7664 197970 7676
rect 295334 7664 295340 7676
rect 197964 7636 295340 7664
rect 197964 7624 197970 7636
rect 295334 7624 295340 7636
rect 295392 7624 295398 7676
rect 347866 7624 347872 7676
rect 347924 7664 347930 7676
rect 367002 7664 367008 7676
rect 347924 7636 367008 7664
rect 347924 7624 347930 7636
rect 367002 7624 367008 7636
rect 367060 7624 367066 7676
rect 176746 7556 176752 7608
rect 176804 7596 176810 7608
rect 288710 7596 288716 7608
rect 176804 7568 288716 7596
rect 176804 7556 176810 7568
rect 288710 7556 288716 7568
rect 288768 7556 288774 7608
rect 310238 7556 310244 7608
rect 310296 7596 310302 7608
rect 329926 7596 329932 7608
rect 310296 7568 329932 7596
rect 310296 7556 310302 7568
rect 329926 7556 329932 7568
rect 329984 7556 329990 7608
rect 347774 7556 347780 7608
rect 347832 7596 347838 7608
rect 369394 7596 369400 7608
rect 347832 7568 369400 7596
rect 347832 7556 347838 7568
rect 369394 7556 369400 7568
rect 369452 7556 369458 7608
rect 380894 7556 380900 7608
rect 380952 7596 380958 7608
rect 476942 7596 476948 7608
rect 380952 7568 476948 7596
rect 380952 7556 380958 7568
rect 476942 7556 476948 7568
rect 477000 7556 477006 7608
rect 3510 6468 3516 6520
rect 3568 6508 3574 6520
rect 8938 6508 8944 6520
rect 3568 6480 8944 6508
rect 3568 6468 3574 6480
rect 8938 6468 8944 6480
rect 8996 6468 9002 6520
rect 367186 6468 367192 6520
rect 367244 6508 367250 6520
rect 430850 6508 430856 6520
rect 367244 6480 430856 6508
rect 367244 6468 367250 6480
rect 430850 6468 430856 6480
rect 430908 6468 430914 6520
rect 368658 6400 368664 6452
rect 368716 6440 368722 6452
rect 434438 6440 434444 6452
rect 368716 6412 434444 6440
rect 368716 6400 368722 6412
rect 434438 6400 434444 6412
rect 434496 6400 434502 6452
rect 369946 6332 369952 6384
rect 370004 6372 370010 6384
rect 437934 6372 437940 6384
rect 370004 6344 437940 6372
rect 370004 6332 370010 6344
rect 437934 6332 437940 6344
rect 437992 6332 437998 6384
rect 235810 6264 235816 6316
rect 235868 6304 235874 6316
rect 306558 6304 306564 6316
rect 235868 6276 306564 6304
rect 235868 6264 235874 6276
rect 306558 6264 306564 6276
rect 306616 6264 306622 6316
rect 371326 6264 371332 6316
rect 371384 6304 371390 6316
rect 441522 6304 441528 6316
rect 371384 6276 441528 6304
rect 371384 6264 371390 6276
rect 441522 6264 441528 6276
rect 441580 6264 441586 6316
rect 237006 6196 237012 6248
rect 237064 6236 237070 6248
rect 304258 6236 304264 6248
rect 237064 6208 304264 6236
rect 237064 6196 237070 6208
rect 304258 6196 304264 6208
rect 304316 6196 304322 6248
rect 345014 6196 345020 6248
rect 345072 6236 345078 6248
rect 359918 6236 359924 6248
rect 345072 6208 359924 6236
rect 345072 6196 345078 6208
rect 359918 6196 359924 6208
rect 359976 6196 359982 6248
rect 371418 6196 371424 6248
rect 371476 6236 371482 6248
rect 445018 6236 445024 6248
rect 371476 6208 445024 6236
rect 371476 6196 371482 6208
rect 445018 6196 445024 6208
rect 445076 6196 445082 6248
rect 128170 6128 128176 6180
rect 128228 6168 128234 6180
rect 231118 6168 231124 6180
rect 128228 6140 231124 6168
rect 128228 6128 128234 6140
rect 231118 6128 231124 6140
rect 231176 6128 231182 6180
rect 306742 6128 306748 6180
rect 306800 6168 306806 6180
rect 328638 6168 328644 6180
rect 306800 6140 328644 6168
rect 306800 6128 306806 6140
rect 328638 6128 328644 6140
rect 328696 6128 328702 6180
rect 346486 6128 346492 6180
rect 346544 6168 346550 6180
rect 364610 6168 364616 6180
rect 346544 6140 364616 6168
rect 346544 6128 346550 6140
rect 364610 6128 364616 6140
rect 364668 6128 364674 6180
rect 412634 6128 412640 6180
rect 412692 6168 412698 6180
rect 576302 6168 576308 6180
rect 412692 6140 576308 6168
rect 412692 6128 412698 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 366358 5516 366364 5568
rect 366416 5556 366422 5568
rect 368198 5556 368204 5568
rect 366416 5528 368204 5556
rect 366416 5516 366422 5528
rect 368198 5516 368204 5528
rect 368256 5516 368262 5568
rect 303154 5040 303160 5092
rect 303212 5080 303218 5092
rect 328546 5080 328552 5092
rect 303212 5052 328552 5080
rect 303212 5040 303218 5052
rect 328546 5040 328552 5052
rect 328604 5040 328610 5092
rect 299658 4972 299664 5024
rect 299716 5012 299722 5024
rect 327258 5012 327264 5024
rect 299716 4984 327264 5012
rect 299716 4972 299722 4984
rect 327258 4972 327264 4984
rect 327316 4972 327322 5024
rect 296070 4904 296076 4956
rect 296128 4944 296134 4956
rect 325786 4944 325792 4956
rect 296128 4916 325792 4944
rect 296128 4904 296134 4916
rect 325786 4904 325792 4916
rect 325844 4904 325850 4956
rect 351178 4904 351184 4956
rect 351236 4944 351242 4956
rect 356330 4944 356336 4956
rect 351236 4916 356336 4944
rect 351236 4904 351242 4916
rect 356330 4904 356336 4916
rect 356388 4904 356394 4956
rect 278314 4836 278320 4888
rect 278372 4876 278378 4888
rect 320358 4876 320364 4888
rect 278372 4848 320364 4876
rect 278372 4836 278378 4848
rect 320358 4836 320364 4848
rect 320416 4836 320422 4888
rect 353294 4836 353300 4888
rect 353352 4876 353358 4888
rect 383562 4876 383568 4888
rect 353352 4848 383568 4876
rect 353352 4836 353358 4848
rect 383562 4836 383568 4848
rect 383620 4836 383626 4888
rect 218146 4768 218152 4820
rect 218204 4808 218210 4820
rect 228358 4808 228364 4820
rect 218204 4780 228364 4808
rect 218204 4768 218210 4780
rect 228358 4768 228364 4780
rect 228416 4768 228422 4820
rect 246390 4768 246396 4820
rect 246448 4808 246454 4820
rect 289078 4808 289084 4820
rect 246448 4780 289084 4808
rect 246448 4768 246454 4780
rect 289078 4768 289084 4780
rect 289136 4768 289142 4820
rect 292574 4768 292580 4820
rect 292632 4808 292638 4820
rect 324498 4808 324504 4820
rect 292632 4780 324504 4808
rect 292632 4768 292638 4780
rect 324498 4768 324504 4780
rect 324556 4768 324562 4820
rect 354674 4768 354680 4820
rect 354732 4808 354738 4820
rect 391842 4808 391848 4820
rect 354732 4780 391848 4808
rect 354732 4768 354738 4780
rect 391842 4768 391848 4780
rect 391900 4768 391906 4820
rect 401594 4768 401600 4820
rect 401652 4808 401658 4820
rect 540790 4808 540796 4820
rect 401652 4780 540796 4808
rect 401652 4768 401658 4780
rect 540790 4768 540796 4780
rect 540848 4768 540854 4820
rect 382918 4496 382924 4548
rect 382976 4536 382982 4548
rect 384758 4536 384764 4548
rect 382976 4508 384764 4536
rect 382976 4496 382982 4508
rect 384758 4496 384764 4508
rect 384816 4496 384822 4548
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 176654 4156 176660 4208
rect 176712 4196 176718 4208
rect 177850 4196 177856 4208
rect 176712 4168 177856 4196
rect 176712 4156 176718 4168
rect 177850 4156 177856 4168
rect 177908 4156 177914 4208
rect 345658 4156 345664 4208
rect 345716 4196 345722 4208
rect 352834 4196 352840 4208
rect 345716 4168 352840 4196
rect 345716 4156 345722 4168
rect 352834 4156 352840 4168
rect 352892 4156 352898 4208
rect 46658 4088 46664 4140
rect 46716 4128 46722 4140
rect 248690 4128 248696 4140
rect 46716 4100 248696 4128
rect 46716 4088 46722 4100
rect 248690 4088 248696 4100
rect 248748 4088 248754 4140
rect 305546 4088 305552 4140
rect 305604 4128 305610 4140
rect 328454 4128 328460 4140
rect 305604 4100 328460 4128
rect 305604 4088 305610 4100
rect 328454 4088 328460 4100
rect 328512 4088 328518 4140
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 336918 4128 336924 4140
rect 332744 4100 336924 4128
rect 332744 4088 332750 4100
rect 336918 4088 336924 4100
rect 336976 4088 336982 4140
rect 341150 4088 341156 4140
rect 341208 4128 341214 4140
rect 345750 4128 345756 4140
rect 341208 4100 345756 4128
rect 341208 4088 341214 4100
rect 345750 4088 345756 4100
rect 345808 4088 345814 4140
rect 367094 4088 367100 4140
rect 367152 4128 367158 4140
rect 429654 4128 429660 4140
rect 367152 4100 429660 4128
rect 367152 4088 367158 4100
rect 429654 4088 429660 4100
rect 429712 4088 429718 4140
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 247310 4060 247316 4072
rect 43128 4032 247316 4060
rect 43128 4020 43134 4032
rect 247310 4020 247316 4032
rect 247368 4020 247374 4072
rect 301958 4020 301964 4072
rect 302016 4060 302022 4072
rect 327074 4060 327080 4072
rect 302016 4032 327080 4060
rect 302016 4020 302022 4032
rect 327074 4020 327080 4032
rect 327132 4020 327138 4072
rect 335538 4060 335544 4072
rect 327276 4032 335544 4060
rect 39574 3952 39580 4004
rect 39632 3992 39638 4004
rect 247126 3992 247132 4004
rect 39632 3964 247132 3992
rect 39632 3952 39638 3964
rect 247126 3952 247132 3964
rect 247184 3952 247190 4004
rect 298462 3952 298468 4004
rect 298520 3992 298526 4004
rect 327166 3992 327172 4004
rect 298520 3964 327172 3992
rect 298520 3952 298526 3964
rect 327166 3952 327172 3964
rect 327224 3952 327230 4004
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 7650 3924 7656 3936
rect 2924 3896 7656 3924
rect 2924 3884 2930 3896
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 35986 3884 35992 3936
rect 36044 3924 36050 3936
rect 245930 3924 245936 3936
rect 36044 3896 245936 3924
rect 36044 3884 36050 3896
rect 245930 3884 245936 3896
rect 245988 3884 245994 3936
rect 294874 3884 294880 3936
rect 294932 3924 294938 3936
rect 325878 3924 325884 3936
rect 294932 3896 325884 3924
rect 294932 3884 294938 3896
rect 325878 3884 325884 3896
rect 325936 3884 325942 3936
rect 326798 3884 326804 3936
rect 326856 3924 326862 3936
rect 327276 3924 327304 4032
rect 335538 4020 335544 4032
rect 335596 4020 335602 4072
rect 340966 4020 340972 4072
rect 341024 4060 341030 4072
rect 346946 4060 346952 4072
rect 341024 4032 346952 4060
rect 341024 4020 341030 4032
rect 346946 4020 346952 4032
rect 347004 4020 347010 4072
rect 368566 4020 368572 4072
rect 368624 4060 368630 4072
rect 433242 4060 433248 4072
rect 368624 4032 433248 4060
rect 368624 4020 368630 4032
rect 433242 4020 433248 4032
rect 433300 4020 433306 4072
rect 333882 3952 333888 4004
rect 333940 3992 333946 4004
rect 337102 3992 337108 4004
rect 333940 3964 337108 3992
rect 333940 3952 333946 3964
rect 337102 3952 337108 3964
rect 337160 3952 337166 4004
rect 368474 3952 368480 4004
rect 368532 3992 368538 4004
rect 436738 3992 436744 4004
rect 368532 3964 436744 3992
rect 368532 3952 368538 3964
rect 436738 3952 436744 3964
rect 436796 3952 436802 4004
rect 326856 3896 327304 3924
rect 326856 3884 326862 3896
rect 327994 3884 328000 3936
rect 328052 3924 328058 3936
rect 335354 3924 335360 3936
rect 328052 3896 335360 3924
rect 328052 3884 328058 3896
rect 335354 3884 335360 3896
rect 335412 3884 335418 3936
rect 342530 3884 342536 3936
rect 342588 3924 342594 3936
rect 348050 3924 348056 3936
rect 342588 3896 348056 3924
rect 342588 3884 342594 3896
rect 348050 3884 348056 3896
rect 348108 3884 348114 3936
rect 369854 3884 369860 3936
rect 369912 3924 369918 3936
rect 440326 3924 440332 3936
rect 369912 3896 440332 3924
rect 369912 3884 369918 3896
rect 440326 3884 440332 3896
rect 440384 3884 440390 3936
rect 32398 3816 32404 3868
rect 32456 3856 32462 3868
rect 244274 3856 244280 3868
rect 32456 3828 244280 3856
rect 32456 3816 32462 3828
rect 244274 3816 244280 3828
rect 244332 3816 244338 3868
rect 291378 3816 291384 3868
rect 291436 3856 291442 3868
rect 324406 3856 324412 3868
rect 291436 3828 324412 3856
rect 291436 3816 291442 3828
rect 324406 3816 324412 3828
rect 324464 3816 324470 3868
rect 329190 3816 329196 3868
rect 329248 3856 329254 3868
rect 335630 3856 335636 3868
rect 329248 3828 335636 3856
rect 329248 3816 329254 3828
rect 335630 3816 335636 3828
rect 335688 3816 335694 3868
rect 342622 3816 342628 3868
rect 342680 3856 342686 3868
rect 350442 3856 350448 3868
rect 342680 3828 350448 3856
rect 342680 3816 342686 3828
rect 350442 3816 350448 3828
rect 350500 3816 350506 3868
rect 371234 3816 371240 3868
rect 371292 3856 371298 3868
rect 443822 3856 443828 3868
rect 371292 3828 443828 3856
rect 371292 3816 371298 3828
rect 443822 3816 443828 3828
rect 443880 3816 443886 3868
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 242894 3788 242900 3800
rect 28960 3760 242900 3788
rect 28960 3748 28966 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 287790 3748 287796 3800
rect 287848 3788 287854 3800
rect 322934 3788 322940 3800
rect 287848 3760 322940 3788
rect 287848 3748 287854 3760
rect 322934 3748 322940 3760
rect 322992 3748 322998 3800
rect 325602 3748 325608 3800
rect 325660 3788 325666 3800
rect 335446 3788 335452 3800
rect 325660 3760 335452 3788
rect 325660 3748 325666 3760
rect 335446 3748 335452 3760
rect 335504 3748 335510 3800
rect 374178 3748 374184 3800
rect 374236 3788 374242 3800
rect 450906 3788 450912 3800
rect 374236 3760 450912 3788
rect 374236 3748 374242 3760
rect 450906 3748 450912 3760
rect 450964 3748 450970 3800
rect 576118 3748 576124 3800
rect 576176 3788 576182 3800
rect 578602 3788 578608 3800
rect 576176 3760 578608 3788
rect 576176 3748 576182 3760
rect 578602 3748 578608 3760
rect 578660 3748 578666 3800
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 24118 3720 24124 3732
rect 14792 3692 24124 3720
rect 14792 3680 14798 3692
rect 24118 3680 24124 3692
rect 24176 3680 24182 3732
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 241514 3720 241520 3732
rect 25372 3692 241520 3720
rect 25372 3680 25378 3692
rect 241514 3680 241520 3692
rect 241572 3680 241578 3732
rect 284294 3680 284300 3732
rect 284352 3720 284358 3732
rect 321554 3720 321560 3732
rect 284352 3692 321560 3720
rect 284352 3680 284358 3692
rect 321554 3680 321560 3692
rect 321612 3680 321618 3732
rect 323302 3680 323308 3732
rect 323360 3720 323366 3732
rect 334158 3720 334164 3732
rect 323360 3692 334164 3720
rect 323360 3680 323366 3692
rect 334158 3680 334164 3692
rect 334216 3680 334222 3732
rect 342438 3680 342444 3732
rect 342496 3720 342502 3732
rect 349246 3720 349252 3732
rect 342496 3692 349252 3720
rect 342496 3680 342502 3692
rect 349246 3680 349252 3692
rect 349304 3680 349310 3732
rect 375374 3680 375380 3732
rect 375432 3720 375438 3732
rect 458082 3720 458088 3732
rect 375432 3692 458088 3720
rect 375432 3680 375438 3692
rect 458082 3680 458088 3692
rect 458140 3680 458146 3732
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 13078 3652 13084 3664
rect 8812 3624 13084 3652
rect 8812 3612 8818 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 241606 3652 241612 3664
rect 24268 3624 241612 3652
rect 24268 3612 24274 3624
rect 241606 3612 241612 3624
rect 241664 3612 241670 3664
rect 280706 3612 280712 3664
rect 280764 3652 280770 3664
rect 321646 3652 321652 3664
rect 280764 3624 321652 3652
rect 280764 3612 280770 3624
rect 321646 3612 321652 3624
rect 321704 3612 321710 3664
rect 322106 3612 322112 3664
rect 322164 3652 322170 3664
rect 334066 3652 334072 3664
rect 322164 3624 334072 3652
rect 322164 3612 322170 3624
rect 334066 3612 334072 3624
rect 334124 3612 334130 3664
rect 346394 3612 346400 3664
rect 346452 3652 346458 3664
rect 362310 3652 362316 3664
rect 346452 3624 362316 3652
rect 346452 3612 346458 3624
rect 362310 3612 362316 3624
rect 362368 3612 362374 3664
rect 378134 3612 378140 3664
rect 378192 3652 378198 3664
rect 465166 3652 465172 3664
rect 378192 3624 465172 3652
rect 378192 3612 378198 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 10318 3584 10324 3596
rect 6512 3556 10324 3584
rect 6512 3544 6518 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 240226 3584 240232 3596
rect 19484 3556 240232 3584
rect 19484 3544 19490 3556
rect 240226 3544 240232 3556
rect 240284 3544 240290 3596
rect 242894 3544 242900 3596
rect 242952 3584 242958 3596
rect 243078 3584 243084 3596
rect 242952 3556 243084 3584
rect 242952 3544 242958 3556
rect 243078 3544 243084 3556
rect 243136 3544 243142 3596
rect 251266 3544 251272 3596
rect 251324 3584 251330 3596
rect 252370 3584 252376 3596
rect 251324 3556 252376 3584
rect 251324 3544 251330 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 273622 3544 273628 3596
rect 273680 3584 273686 3596
rect 318794 3584 318800 3596
rect 273680 3556 318800 3584
rect 273680 3544 273686 3556
rect 318794 3544 318800 3556
rect 318852 3544 318858 3596
rect 319714 3544 319720 3596
rect 319772 3584 319778 3596
rect 332594 3584 332600 3596
rect 319772 3556 332600 3584
rect 319772 3544 319778 3556
rect 332594 3544 332600 3556
rect 332652 3544 332658 3596
rect 342346 3544 342352 3596
rect 342404 3584 342410 3596
rect 351638 3584 351644 3596
rect 342404 3556 351644 3584
rect 342404 3544 342410 3556
rect 351638 3544 351644 3556
rect 351696 3544 351702 3596
rect 360194 3544 360200 3596
rect 360252 3584 360258 3596
rect 408402 3584 408408 3596
rect 360252 3556 408408 3584
rect 360252 3544 360258 3556
rect 408402 3544 408408 3556
rect 408460 3544 408466 3596
rect 414198 3544 414204 3596
rect 414256 3584 414262 3596
rect 582190 3584 582196 3596
rect 414256 3556 582196 3584
rect 414256 3544 414262 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 3418 3516 3424 3528
rect 624 3488 3424 3516
rect 624 3476 630 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 15838 3516 15844 3528
rect 12400 3488 15844 3516
rect 12400 3476 12406 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 240410 3516 240416 3528
rect 20680 3488 240416 3516
rect 20680 3476 20686 3488
rect 240410 3476 240416 3488
rect 240468 3476 240474 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 316310 3516 316316 3528
rect 266596 3488 316316 3516
rect 266596 3476 266602 3488
rect 316310 3476 316316 3488
rect 316368 3476 316374 3528
rect 318518 3476 318524 3528
rect 318576 3516 318582 3528
rect 332502 3516 332508 3528
rect 318576 3488 332508 3516
rect 318576 3476 318582 3488
rect 332502 3476 332508 3488
rect 332560 3476 332566 3528
rect 337470 3476 337476 3528
rect 337528 3516 337534 3528
rect 338390 3516 338396 3528
rect 337528 3488 338396 3516
rect 337528 3476 337534 3488
rect 338390 3476 338396 3488
rect 338448 3476 338454 3528
rect 338666 3476 338672 3528
rect 338724 3516 338730 3528
rect 339586 3516 339592 3528
rect 338724 3488 339592 3516
rect 338724 3476 338730 3488
rect 339586 3476 339592 3488
rect 339644 3476 339650 3528
rect 339678 3476 339684 3528
rect 339736 3516 339742 3528
rect 340966 3516 340972 3528
rect 339736 3488 340972 3516
rect 339736 3476 339742 3488
rect 340966 3476 340972 3488
rect 341024 3476 341030 3528
rect 343726 3476 343732 3528
rect 343784 3516 343790 3528
rect 354030 3516 354036 3528
rect 343784 3488 354036 3516
rect 343784 3476 343790 3488
rect 354030 3476 354036 3488
rect 354088 3476 354094 3528
rect 357434 3476 357440 3528
rect 357492 3516 357498 3528
rect 358722 3516 358728 3528
rect 357492 3488 358728 3516
rect 357492 3476 357498 3488
rect 358722 3476 358728 3488
rect 358780 3476 358786 3528
rect 373994 3476 374000 3528
rect 374052 3516 374058 3528
rect 375282 3516 375288 3528
rect 374052 3488 375288 3516
rect 374052 3476 374058 3488
rect 375282 3476 375288 3488
rect 375340 3476 375346 3528
rect 379514 3476 379520 3528
rect 379572 3516 379578 3528
rect 472250 3516 472256 3528
rect 379572 3488 472256 3516
rect 379572 3476 379578 3488
rect 472250 3476 472256 3488
rect 472308 3476 472314 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 4798 3448 4804 3460
rect 1728 3420 4804 3448
rect 1728 3408 1734 3420
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 14550 3448 14556 3460
rect 10008 3420 14556 3448
rect 10008 3408 10014 3420
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 238754 3448 238760 3460
rect 15988 3420 238760 3448
rect 15988 3408 15994 3420
rect 238754 3408 238760 3420
rect 238812 3408 238818 3460
rect 299474 3408 299480 3460
rect 299532 3448 299538 3460
rect 300762 3448 300768 3460
rect 299532 3420 300768 3448
rect 299532 3408 299538 3420
rect 300762 3408 300768 3420
rect 300820 3408 300826 3460
rect 316218 3408 316224 3460
rect 316276 3448 316282 3460
rect 331490 3448 331496 3460
rect 316276 3420 331496 3448
rect 316276 3408 316282 3420
rect 331490 3408 331496 3420
rect 331548 3408 331554 3460
rect 343634 3408 343640 3460
rect 343692 3448 343698 3460
rect 355226 3448 355232 3460
rect 343692 3420 355232 3448
rect 343692 3408 343698 3420
rect 355226 3408 355232 3420
rect 355284 3408 355290 3460
rect 361574 3408 361580 3460
rect 361632 3448 361638 3460
rect 411898 3448 411904 3460
rect 361632 3420 411904 3448
rect 361632 3408 361638 3420
rect 411898 3408 411904 3420
rect 411956 3408 411962 3460
rect 415394 3408 415400 3460
rect 415452 3448 415458 3460
rect 416682 3448 416688 3460
rect 415452 3420 416688 3448
rect 415452 3408 415458 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 416774 3408 416780 3460
rect 416832 3448 416838 3460
rect 580994 3448 581000 3460
rect 416832 3420 581000 3448
rect 416832 3408 416838 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 77294 3340 77300 3392
rect 77352 3380 77358 3392
rect 78214 3380 78220 3392
rect 77352 3352 78220 3380
rect 77352 3340 77358 3352
rect 78214 3340 78220 3352
rect 78272 3340 78278 3392
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 269114 3380 269120 3392
rect 120000 3352 269120 3380
rect 7650 3272 7656 3324
rect 7708 3312 7714 3324
rect 11698 3312 11704 3324
rect 7708 3284 11704 3312
rect 7708 3272 7714 3284
rect 11698 3272 11704 3284
rect 11756 3272 11762 3324
rect 114002 3272 114008 3324
rect 114060 3312 114066 3324
rect 120000 3312 120028 3352
rect 269114 3340 269120 3352
rect 269172 3340 269178 3392
rect 309042 3340 309048 3392
rect 309100 3380 309106 3392
rect 329834 3380 329840 3392
rect 309100 3352 329840 3380
rect 309100 3340 309106 3352
rect 329834 3340 329840 3352
rect 329892 3340 329898 3392
rect 341058 3340 341064 3392
rect 341116 3380 341122 3392
rect 344554 3380 344560 3392
rect 341116 3352 344560 3380
rect 341116 3340 341122 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 426158 3380 426164 3392
rect 365772 3352 426164 3380
rect 365772 3340 365778 3352
rect 426158 3340 426164 3352
rect 426216 3340 426222 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 114060 3284 120028 3312
rect 114060 3272 114066 3284
rect 121086 3272 121092 3324
rect 121144 3312 121150 3324
rect 272150 3312 272156 3324
rect 121144 3284 272156 3312
rect 121144 3272 121150 3284
rect 272150 3272 272156 3284
rect 272208 3272 272214 3324
rect 312630 3272 312636 3324
rect 312688 3312 312694 3324
rect 331306 3312 331312 3324
rect 312688 3284 331312 3312
rect 312688 3272 312694 3284
rect 331306 3272 331312 3284
rect 331364 3272 331370 3324
rect 364426 3272 364432 3324
rect 364484 3312 364490 3324
rect 422570 3312 422576 3324
rect 364484 3284 422576 3312
rect 364484 3272 364490 3284
rect 422570 3272 422576 3284
rect 422628 3272 422634 3324
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 273438 3244 273444 3256
rect 124732 3216 273444 3244
rect 124732 3204 124738 3216
rect 273438 3204 273444 3216
rect 273496 3204 273502 3256
rect 315022 3204 315028 3256
rect 315080 3244 315086 3256
rect 331398 3244 331404 3256
rect 315080 3216 331404 3244
rect 315080 3204 315086 3216
rect 331398 3204 331404 3216
rect 331456 3204 331462 3256
rect 336826 3244 336832 3256
rect 335326 3216 336832 3244
rect 218054 3136 218060 3188
rect 218112 3176 218118 3188
rect 219250 3176 219256 3188
rect 218112 3148 219256 3176
rect 218112 3136 218118 3148
rect 219250 3136 219256 3148
rect 219308 3136 219314 3188
rect 270034 3136 270040 3188
rect 270092 3176 270098 3188
rect 317690 3176 317696 3188
rect 270092 3148 317696 3176
rect 270092 3136 270098 3148
rect 317690 3136 317696 3148
rect 317748 3136 317754 3188
rect 330386 3136 330392 3188
rect 330444 3176 330450 3188
rect 335326 3176 335354 3216
rect 336826 3204 336832 3216
rect 336884 3204 336890 3256
rect 364334 3204 364340 3256
rect 364392 3244 364398 3256
rect 418982 3244 418988 3256
rect 364392 3216 418988 3244
rect 364392 3204 364398 3216
rect 418982 3204 418988 3216
rect 419040 3204 419046 3256
rect 330444 3148 335354 3176
rect 330444 3136 330450 3148
rect 336274 3136 336280 3188
rect 336332 3176 336338 3188
rect 338206 3176 338212 3188
rect 336332 3148 338212 3176
rect 336332 3136 336338 3148
rect 338206 3136 338212 3148
rect 338264 3136 338270 3188
rect 398926 3136 398932 3188
rect 398984 3176 398990 3188
rect 400122 3176 400128 3188
rect 398984 3148 400128 3176
rect 398984 3136 398990 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 414106 3136 414112 3188
rect 414164 3176 414170 3188
rect 416774 3176 416780 3188
rect 414164 3148 416780 3176
rect 414164 3136 414170 3148
rect 416774 3136 416780 3148
rect 416832 3136 416838 3188
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 6270 2904 6276 2916
rect 4120 2876 6276 2904
rect 4120 2864 4126 2876
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 423674 960 423680 1012
rect 423732 1000 423738 1012
rect 424962 1000 424968 1012
rect 423732 972 424968 1000
rect 423732 960 423738 972
rect 424962 960 424968 972
rect 425020 960 425026 1012
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 283840 700816 283892 700868
rect 328460 700816 328512 700868
rect 318800 700748 318852 700800
rect 413652 700748 413704 700800
rect 218980 700680 219032 700732
rect 332600 700680 332652 700732
rect 314660 700612 314712 700664
rect 478512 700612 478564 700664
rect 154120 700544 154172 700596
rect 338120 700544 338172 700596
rect 89168 700476 89220 700528
rect 342260 700476 342312 700528
rect 72976 700408 73028 700460
rect 340880 700408 340932 700460
rect 24308 700340 24360 700392
rect 347872 700340 347924 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 478144 700272 478196 700324
rect 559656 700272 559708 700324
rect 235172 698912 235224 698964
rect 329840 698912 329892 698964
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 303620 696940 303672 696992
rect 580172 696940 580224 696992
rect 305000 683136 305052 683188
rect 580172 683136 580224 683188
rect 300860 670760 300912 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 351920 670692 351972 670744
rect 3516 656888 3568 656940
rect 350540 656888 350592 656940
rect 298100 643084 298152 643136
rect 580172 643084 580224 643136
rect 299572 630640 299624 630692
rect 580172 630640 580224 630692
rect 3332 618264 3384 618316
rect 356060 618264 356112 618316
rect 296720 616836 296772 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 354680 605820 354732 605872
rect 293960 590656 294012 590708
rect 579804 590656 579856 590708
rect 295340 576852 295392 576904
rect 580172 576852 580224 576904
rect 3056 565836 3108 565888
rect 361580 565836 361632 565888
rect 292580 563048 292632 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 360200 553392 360252 553444
rect 288440 536800 288492 536852
rect 580172 536800 580224 536852
rect 289820 524424 289872 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 365720 514768 365772 514820
rect 287060 510620 287112 510672
rect 580172 510620 580224 510672
rect 320180 502936 320232 502988
rect 364340 502936 364392 502988
rect 3240 500964 3292 501016
rect 364340 500964 364392 501016
rect 284300 484372 284352 484424
rect 580172 484372 580224 484424
rect 285864 470568 285916 470620
rect 579988 470568 580040 470620
rect 169760 468460 169812 468512
rect 334808 468460 334860 468512
rect 299480 467100 299532 467152
rect 325700 467100 325752 467152
rect 316040 465672 316092 465724
rect 429200 465672 429252 465724
rect 311164 464312 311216 464364
rect 494060 464312 494112 464364
rect 226984 462476 227036 462528
rect 375932 462476 375984 462528
rect 277124 462408 277176 462460
rect 425704 462408 425756 462460
rect 3516 462340 3568 462392
rect 371240 462340 371292 462392
rect 307116 461592 307168 461644
rect 478144 461592 478196 461644
rect 233976 461320 234028 461372
rect 369860 461320 369912 461372
rect 280068 461252 280120 461304
rect 417516 461252 417568 461304
rect 278688 461184 278740 461236
rect 422944 461184 422996 461236
rect 273996 461116 274048 461168
rect 421564 461116 421616 461168
rect 228364 461048 228416 461100
rect 379152 461048 379204 461100
rect 229744 460980 229796 461032
rect 396540 460980 396592 461032
rect 4896 460912 4948 460964
rect 391940 460912 391992 460964
rect 318156 460844 318208 460896
rect 397460 460844 397512 460896
rect 201500 460776 201552 460828
rect 331772 460776 331824 460828
rect 313096 460708 313148 460760
rect 462320 460708 462372 460760
rect 136640 460640 136692 460692
rect 336740 460640 336792 460692
rect 308680 460572 308732 460624
rect 527180 460572 527232 460624
rect 310244 460504 310296 460556
rect 542360 460504 542412 460556
rect 104900 460436 104952 460488
rect 339684 460436 339736 460488
rect 3608 460368 3660 460420
rect 353852 460368 353904 460420
rect 3700 460300 3752 460352
rect 358820 460300 358872 460352
rect 3792 460232 3844 460284
rect 363328 460232 363380 460284
rect 3884 460164 3936 460216
rect 368112 460164 368164 460216
rect 266360 460096 266412 460148
rect 327080 460096 327132 460148
rect 324136 460028 324188 460080
rect 347780 460028 347832 460080
rect 322848 459960 322900 460012
rect 331220 459960 331272 460012
rect 349804 459620 349856 459672
rect 374368 459620 374420 459672
rect 349068 459552 349120 459604
rect 380900 459552 380952 459604
rect 3424 458804 3476 458856
rect 349068 458804 349120 458856
rect 233884 458736 233936 458788
rect 377588 458736 377640 458788
rect 275560 458668 275612 458720
rect 424324 458668 424376 458720
rect 232504 458600 232556 458652
rect 382280 458600 382332 458652
rect 231216 458532 231268 458584
rect 387064 458532 387116 458584
rect 255044 458464 255096 458516
rect 420184 458464 420236 458516
rect 245568 458396 245620 458448
rect 418804 458396 418856 458448
rect 240784 458328 240836 458380
rect 417424 458328 417476 458380
rect 235908 458260 235960 458312
rect 580264 458260 580316 458312
rect 3608 458192 3660 458244
rect 373126 458192 373178 458244
rect 3516 457444 3568 457496
rect 281632 457580 281684 457632
rect 283380 457444 283432 457496
rect 349804 457444 349856 457496
rect 427084 456832 427136 456884
rect 580172 456764 580224 456816
rect 3332 449828 3384 449880
rect 233976 449828 234028 449880
rect 417516 431876 417568 431928
rect 580172 431876 580224 431928
rect 427084 419432 427136 419484
rect 580172 419432 580224 419484
rect 2964 411204 3016 411256
rect 226984 411204 227036 411256
rect 422944 405628 422996 405680
rect 579620 405628 579672 405680
rect 424324 379448 424376 379500
rect 580172 379448 580224 379500
rect 3516 372512 3568 372564
rect 233884 372512 233936 372564
rect 425704 365644 425756 365696
rect 580172 365644 580224 365696
rect 421564 353200 421616 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 228364 346332 228416 346384
rect 270546 337764 270598 337816
rect 270776 337764 270828 337816
rect 331220 336880 331272 336932
rect 331588 336880 331640 336932
rect 294420 336744 294472 336796
rect 399024 336744 399076 336796
rect 242992 336676 243044 336728
rect 243268 336676 243320 336728
rect 246304 336676 246356 336728
rect 247224 336676 247276 336728
rect 251824 336676 251876 336728
rect 254216 336676 254268 336728
rect 269764 336676 269816 336728
rect 273536 336676 273588 336728
rect 282828 336676 282880 336728
rect 285680 336676 285732 336728
rect 287704 336676 287756 336728
rect 290372 336676 290424 336728
rect 293224 336676 293276 336728
rect 300768 336676 300820 336728
rect 304080 336676 304132 336728
rect 307024 336676 307076 336728
rect 313372 336676 313424 336728
rect 316132 336676 316184 336728
rect 316316 336676 316368 336728
rect 342444 336676 342496 336728
rect 342628 336676 342680 336728
rect 346400 336676 346452 336728
rect 346676 336676 346728 336728
rect 367100 336676 367152 336728
rect 367468 336676 367520 336728
rect 386420 336676 386472 336728
rect 386788 336676 386840 336728
rect 291936 336608 291988 336660
rect 293316 336608 293368 336660
rect 298744 336608 298796 336660
rect 307116 336608 307168 336660
rect 314844 336608 314896 336660
rect 244924 336540 244976 336592
rect 246212 336540 246264 336592
rect 294604 336540 294656 336592
rect 340788 336540 340840 336592
rect 341340 336540 341392 336592
rect 401600 336676 401652 336728
rect 401876 336676 401928 336728
rect 400864 336540 400916 336592
rect 298744 336472 298796 336524
rect 302424 336472 302476 336524
rect 302976 336472 303028 336524
rect 309692 336472 309744 336524
rect 350080 336472 350132 336524
rect 358084 336472 358136 336524
rect 362868 336472 362920 336524
rect 373356 336472 373408 336524
rect 353760 336404 353812 336456
rect 382924 336404 382976 336456
rect 402336 336404 402388 336456
rect 417516 336404 417568 336456
rect 231124 336336 231176 336388
rect 274272 336336 274324 336388
rect 358176 336336 358228 336388
rect 387064 336336 387116 336388
rect 396448 336336 396500 336388
rect 424324 336336 424376 336388
rect 228364 336268 228416 336320
rect 302240 336268 302292 336320
rect 315304 336268 315356 336320
rect 324320 336268 324372 336320
rect 334348 336268 334400 336320
rect 338212 336268 338264 336320
rect 345664 336268 345716 336320
rect 357440 336268 357492 336320
rect 362776 336268 362828 336320
rect 370504 336268 370556 336320
rect 373080 336268 373132 336320
rect 447140 336268 447192 336320
rect 117320 336200 117372 336252
rect 271052 336200 271104 336252
rect 276664 336200 276716 336252
rect 277952 336200 278004 336252
rect 302884 336200 302936 336252
rect 316684 336200 316736 336252
rect 339500 336200 339552 336252
rect 339684 336200 339736 336252
rect 347320 336200 347372 336252
rect 362960 336200 363012 336252
rect 375288 336200 375340 336252
rect 454040 336200 454092 336252
rect 110420 336132 110472 336184
rect 268844 336132 268896 336184
rect 297364 336132 297416 336184
rect 311900 336132 311952 336184
rect 324320 336132 324372 336184
rect 334900 336132 334952 336184
rect 343824 336132 343876 336184
rect 345664 336132 345716 336184
rect 348608 336132 348660 336184
rect 366272 336132 366324 336184
rect 377220 336132 377272 336184
rect 460940 336132 460992 336184
rect 102140 336064 102192 336116
rect 10324 335996 10376 336048
rect 236644 335996 236696 336048
rect 264244 336064 264296 336116
rect 264980 336064 265032 336116
rect 289084 336064 289136 336116
rect 310796 336064 310848 336116
rect 318064 336064 318116 336116
rect 331220 336064 331272 336116
rect 350816 336064 350868 336116
rect 374000 336064 374052 336116
rect 379888 336064 379940 336116
rect 467840 336064 467892 336116
rect 266728 335996 266780 336048
rect 276756 335996 276808 336048
rect 284484 335996 284536 336048
rect 286232 335996 286284 336048
rect 291200 335996 291252 336048
rect 291844 335996 291896 336048
rect 315212 335996 315264 336048
rect 320180 335996 320232 336048
rect 333980 335996 334032 336048
rect 344928 335996 344980 336048
rect 351184 335996 351236 336048
rect 351920 335996 351972 336048
rect 377404 335996 377456 336048
rect 381820 335996 381872 336048
rect 474740 335996 474792 336048
rect 260840 335928 260892 335980
rect 261116 335928 261168 335980
rect 305644 335928 305696 335980
rect 307208 335928 307260 335980
rect 271144 335792 271196 335844
rect 272432 335792 272484 335844
rect 319444 335792 319496 335844
rect 321008 335792 321060 335844
rect 286416 335724 286468 335776
rect 287796 335724 287848 335776
rect 320824 335724 320876 335776
rect 326528 335724 326580 335776
rect 297456 335656 297508 335708
rect 299848 335656 299900 335708
rect 340972 335656 341024 335708
rect 342260 335656 342312 335708
rect 303528 335588 303580 335640
rect 306472 335588 306524 335640
rect 289176 335520 289228 335572
rect 290004 335520 290056 335572
rect 411812 335452 411864 335504
rect 413284 335452 413336 335504
rect 301504 335384 301556 335436
rect 308588 335384 308640 335436
rect 379980 335384 380032 335436
rect 381544 335384 381596 335436
rect 233976 335316 234028 335368
rect 240140 335316 240192 335368
rect 295984 335316 296036 335368
rect 296720 335316 296772 335368
rect 304264 335316 304316 335368
rect 307852 335316 307904 335368
rect 313924 335316 313976 335368
rect 317420 335316 317472 335368
rect 331588 335316 331640 335368
rect 337108 335316 337160 335368
rect 224960 334636 225012 334688
rect 300768 334636 300820 334688
rect 383568 334636 383620 334688
rect 480260 334636 480312 334688
rect 3424 334568 3476 334620
rect 234804 334568 234856 334620
rect 405280 334568 405332 334620
rect 550640 334568 550692 334620
rect 384488 333276 384540 333328
rect 483020 333276 483072 333328
rect 231860 333140 231912 333192
rect 303528 333208 303580 333260
rect 408592 333140 408644 333192
rect 561680 333208 561732 333260
rect 175280 331916 175332 331968
rect 288900 331916 288952 331968
rect 46940 331848 46992 331900
rect 249432 331848 249484 331900
rect 397552 331848 397604 331900
rect 525800 331848 525852 331900
rect 280436 331168 280488 331220
rect 280620 331168 280672 331220
rect 283196 330760 283248 330812
rect 283472 330760 283524 330812
rect 168380 330556 168432 330608
rect 57980 330488 58032 330540
rect 252744 330624 252796 330676
rect 286692 330556 286744 330608
rect 390008 330556 390060 330608
rect 500960 330556 501012 330608
rect 249800 330488 249852 330540
rect 250168 330488 250220 330540
rect 251180 330488 251232 330540
rect 252008 330488 252060 330540
rect 254032 330488 254084 330540
rect 254952 330488 255004 330540
rect 255412 330488 255464 330540
rect 255688 330488 255740 330540
rect 256700 330488 256752 330540
rect 257160 330488 257212 330540
rect 258172 330488 258224 330540
rect 258632 330488 258684 330540
rect 260932 330488 260984 330540
rect 261852 330488 261904 330540
rect 262312 330488 262364 330540
rect 263324 330488 263376 330540
rect 266544 330488 266596 330540
rect 267004 330488 267056 330540
rect 267832 330488 267884 330540
rect 268476 330488 268528 330540
rect 269120 330488 269172 330540
rect 269948 330488 270000 330540
rect 270592 330488 270644 330540
rect 271328 330488 271380 330540
rect 271972 330488 272024 330540
rect 272800 330488 272852 330540
rect 285772 330488 285824 330540
rect 286324 330488 286376 330540
rect 287152 330488 287204 330540
rect 288164 330488 288216 330540
rect 291384 330488 291436 330540
rect 292212 330488 292264 330540
rect 294236 330488 294288 330540
rect 295156 330488 295208 330540
rect 295340 330488 295392 330540
rect 295800 330488 295852 330540
rect 298376 330488 298428 330540
rect 299112 330488 299164 330540
rect 299572 330488 299624 330540
rect 300584 330488 300636 330540
rect 300860 330488 300912 330540
rect 301688 330488 301740 330540
rect 313464 330488 313516 330540
rect 314108 330488 314160 330540
rect 317696 330488 317748 330540
rect 318156 330488 318208 330540
rect 318800 330488 318852 330540
rect 319260 330488 319312 330540
rect 332600 330488 332652 330540
rect 333060 330488 333112 330540
rect 335360 330488 335412 330540
rect 336004 330488 336056 330540
rect 360200 330488 360252 330540
rect 360844 330488 360896 330540
rect 363144 330488 363196 330540
rect 363788 330488 363840 330540
rect 364432 330488 364484 330540
rect 365260 330488 365312 330540
rect 365812 330488 365864 330540
rect 366732 330488 366784 330540
rect 368480 330488 368532 330540
rect 369584 330488 369636 330540
rect 390744 330488 390796 330540
rect 391204 330488 391256 330540
rect 392032 330488 392084 330540
rect 392584 330488 392636 330540
rect 393412 330488 393464 330540
rect 394424 330488 394476 330540
rect 394700 330488 394752 330540
rect 395160 330488 395212 330540
rect 397460 330488 397512 330540
rect 398104 330488 398156 330540
rect 408500 330488 408552 330540
rect 409052 330488 409104 330540
rect 409972 330488 410024 330540
rect 410892 330488 410944 330540
rect 411352 330488 411404 330540
rect 412364 330488 412416 330540
rect 244280 330420 244332 330472
rect 244740 330420 244792 330472
rect 249892 330420 249944 330472
rect 250904 330420 250956 330472
rect 255320 330420 255372 330472
rect 256424 330420 256476 330472
rect 256792 330420 256844 330472
rect 257528 330420 257580 330472
rect 258264 330420 258316 330472
rect 259000 330420 259052 330472
rect 266452 330420 266504 330472
rect 267372 330420 267424 330472
rect 317512 330420 317564 330472
rect 318524 330420 318576 330472
rect 318984 330420 319036 330472
rect 319904 330420 319956 330472
rect 332692 330420 332744 330472
rect 333428 330420 333480 330472
rect 390560 330420 390612 330472
rect 391480 330420 391532 330472
rect 391940 330420 391992 330472
rect 392952 330420 393004 330472
rect 410432 330420 410484 330472
rect 567200 330488 567252 330540
rect 258080 330352 258132 330404
rect 258448 330352 258500 330404
rect 296996 330352 297048 330404
rect 297640 330352 297692 330404
rect 361580 329672 361632 329724
rect 361948 329672 362000 329724
rect 396172 329672 396224 329724
rect 397000 329672 397052 329724
rect 262220 329264 262272 329316
rect 262956 329264 263008 329316
rect 164240 329128 164292 329180
rect 282828 329128 282880 329180
rect 283012 329128 283064 329180
rect 283748 329128 283800 329180
rect 60740 329060 60792 329112
rect 253940 329060 253992 329112
rect 367284 329060 367336 329112
rect 368112 329060 368164 329112
rect 392124 329060 392176 329112
rect 507860 329060 507912 329112
rect 314844 328788 314896 328840
rect 315580 328788 315632 328840
rect 295432 328720 295484 328772
rect 296168 328720 296220 328772
rect 245752 328516 245804 328568
rect 246580 328516 246632 328568
rect 265164 327972 265216 328024
rect 265900 327972 265952 328024
rect 365720 327836 365772 327888
rect 366364 327836 366416 327888
rect 201500 327768 201552 327820
rect 296720 327768 296772 327820
rect 396080 327768 396132 327820
rect 396632 327768 396684 327820
rect 125600 327700 125652 327752
rect 269764 327700 269816 327752
rect 394056 327700 394108 327752
rect 514760 327700 514812 327752
rect 259552 327632 259604 327684
rect 260380 327632 260432 327684
rect 367192 327632 367244 327684
rect 367744 327632 367796 327684
rect 393320 327632 393372 327684
rect 393688 327632 393740 327684
rect 378324 326680 378376 326732
rect 383752 326680 383804 326732
rect 237564 326476 237616 326528
rect 237748 326476 237800 326528
rect 241796 326476 241848 326528
rect 241980 326476 242032 326528
rect 354956 326476 355008 326528
rect 355140 326476 355192 326528
rect 375564 326476 375616 326528
rect 375748 326476 375800 326528
rect 378324 326476 378376 326528
rect 381084 326476 381136 326528
rect 381268 326476 381320 326528
rect 383844 326476 383896 326528
rect 193220 326408 193272 326460
rect 293224 326408 293276 326460
rect 323032 326408 323084 326460
rect 323952 326408 324004 326460
rect 328460 326408 328512 326460
rect 329104 326408 329156 326460
rect 329932 326408 329984 326460
rect 330576 326408 330628 326460
rect 354680 326408 354732 326460
rect 355692 326408 355744 326460
rect 356244 326408 356296 326460
rect 356428 326408 356480 326460
rect 369860 326408 369912 326460
rect 370688 326408 370740 326460
rect 371424 326408 371476 326460
rect 372160 326408 372212 326460
rect 372712 326408 372764 326460
rect 373632 326408 373684 326460
rect 374184 326408 374236 326460
rect 374736 326408 374788 326460
rect 375380 326408 375432 326460
rect 376208 326408 376260 326460
rect 376852 326408 376904 326460
rect 377036 326408 377088 326460
rect 379520 326408 379572 326460
rect 380532 326408 380584 326460
rect 380900 326408 380952 326460
rect 382004 326408 382056 326460
rect 383752 326408 383804 326460
rect 384580 326408 384632 326460
rect 385224 326408 385276 326460
rect 385684 326408 385736 326460
rect 386604 326408 386656 326460
rect 387524 326408 387576 326460
rect 387892 326408 387944 326460
rect 388260 326408 388312 326460
rect 401692 326408 401744 326460
rect 402520 326408 402572 326460
rect 403072 326408 403124 326460
rect 403532 326408 403584 326460
rect 404452 326408 404504 326460
rect 404636 326408 404688 326460
rect 405924 326408 405976 326460
rect 406476 326408 406528 326460
rect 407120 326408 407172 326460
rect 407580 326408 407632 326460
rect 11704 326340 11756 326392
rect 237012 326340 237064 326392
rect 237380 326340 237432 326392
rect 238116 326340 238168 326392
rect 238760 326340 238812 326392
rect 239588 326340 239640 326392
rect 240232 326340 240284 326392
rect 240692 326340 240744 326392
rect 241612 326340 241664 326392
rect 242164 326340 242216 326392
rect 274640 326340 274692 326392
rect 275008 326340 275060 326392
rect 276020 326340 276072 326392
rect 276480 326340 276532 326392
rect 277492 326340 277544 326392
rect 278320 326340 278372 326392
rect 278964 326340 279016 326392
rect 279424 326340 279476 326392
rect 280344 326340 280396 326392
rect 281264 326340 281316 326392
rect 281540 326340 281592 326392
rect 282000 326340 282052 326392
rect 305000 326340 305052 326392
rect 306104 326340 306156 326392
rect 306564 326340 306616 326392
rect 307484 326340 307536 326392
rect 309324 326340 309376 326392
rect 310060 326340 310112 326392
rect 310612 326340 310664 326392
rect 311164 326340 311216 326392
rect 321560 326340 321612 326392
rect 322480 326340 322532 326392
rect 322940 326340 322992 326392
rect 323584 326340 323636 326392
rect 327080 326340 327132 326392
rect 328000 326340 328052 326392
rect 328644 326340 328696 326392
rect 329472 326340 329524 326392
rect 329840 326340 329892 326392
rect 330208 326340 330260 326392
rect 340972 326340 341024 326392
rect 341892 326340 341944 326392
rect 342352 326340 342404 326392
rect 343272 326340 343324 326392
rect 346492 326340 346544 326392
rect 347412 326340 347464 326392
rect 350540 326340 350592 326392
rect 351368 326340 351420 326392
rect 354772 326340 354824 326392
rect 355324 326340 355376 326392
rect 356060 326340 356112 326392
rect 357164 326340 357216 326392
rect 357532 326340 357584 326392
rect 358268 326340 358320 326392
rect 364616 326340 364668 326392
rect 419540 326340 419592 326392
rect 241520 326272 241572 326324
rect 242532 326272 242584 326324
rect 278780 326272 278832 326324
rect 279792 326272 279844 326324
rect 280160 326272 280212 326324
rect 280896 326272 280948 326324
rect 371240 326272 371292 326324
rect 371792 326272 371844 326324
rect 378232 326272 378284 326324
rect 379152 326272 379204 326324
rect 387800 326272 387852 326324
rect 388628 326272 388680 326324
rect 402980 326272 403032 326324
rect 403900 326272 403952 326324
rect 405740 326272 405792 326324
rect 406844 326272 406896 326324
rect 407212 326272 407264 326324
rect 407948 326272 408000 326324
rect 242900 326000 242952 326052
rect 243636 326000 243688 326052
rect 176660 324980 176712 325032
rect 289912 324980 289964 325032
rect 160100 324912 160152 324964
rect 276756 324912 276808 324964
rect 365996 324912 366048 324964
rect 423680 324912 423732 324964
rect 292580 324844 292632 324896
rect 292764 324844 292816 324896
rect 347780 323824 347832 323876
rect 348792 323824 348844 323876
rect 386512 323824 386564 323876
rect 387156 323824 387208 323876
rect 385040 323688 385092 323740
rect 386052 323688 386104 323740
rect 128360 323620 128412 323672
rect 274824 323620 274876 323672
rect 26240 323552 26292 323604
rect 243176 323552 243228 323604
rect 305184 323552 305236 323604
rect 305368 323552 305420 323604
rect 358820 323552 358872 323604
rect 359096 323552 359148 323604
rect 378140 323552 378192 323604
rect 378416 323552 378468 323604
rect 398472 323552 398524 323604
rect 529940 323552 529992 323604
rect 302424 323280 302476 323332
rect 303160 323280 303212 323332
rect 343640 323280 343692 323332
rect 344376 323280 344428 323332
rect 358912 323212 358964 323264
rect 359740 323212 359792 323264
rect 305092 322464 305144 322516
rect 305736 322464 305788 322516
rect 403164 322464 403216 322516
rect 403348 322464 403400 322516
rect 189080 322260 189132 322312
rect 291936 322260 291988 322312
rect 51080 322192 51132 322244
rect 250536 322192 250588 322244
rect 345020 322192 345072 322244
rect 345848 322192 345900 322244
rect 398932 322192 398984 322244
rect 532700 322192 532752 322244
rect 273352 322056 273404 322108
rect 273904 322056 273956 322108
rect 347872 321512 347924 321564
rect 348056 321512 348108 321564
rect 367376 320900 367428 320952
rect 427820 320900 427872 320952
rect 215300 320832 215352 320884
rect 301320 320832 301372 320884
rect 385316 320832 385368 320884
rect 487160 320832 487212 320884
rect 248420 320764 248472 320816
rect 248604 320764 248656 320816
rect 3516 320084 3568 320136
rect 232504 320084 232556 320136
rect 325792 319472 325844 319524
rect 325976 319472 326028 319524
rect 369216 319472 369268 319524
rect 434720 319472 434772 319524
rect 205640 319404 205692 319456
rect 298284 319404 298336 319456
rect 386696 319404 386748 319456
rect 489920 319404 489972 319456
rect 371516 318112 371568 318164
rect 441620 318112 441672 318164
rect 219440 318044 219492 318096
rect 302332 318044 302384 318096
rect 386604 318044 386656 318096
rect 494060 318044 494112 318096
rect 223580 316684 223632 316736
rect 303804 316684 303856 316736
rect 387800 316684 387852 316736
rect 498200 316684 498252 316736
rect 226340 315256 226392 315308
rect 305276 315256 305328 315308
rect 394700 315256 394752 315308
rect 518900 315256 518952 315308
rect 118700 313896 118752 313948
rect 272064 313896 272116 313948
rect 391940 313896 391992 313948
rect 512000 313896 512052 313948
rect 171140 312604 171192 312656
rect 286416 312604 286468 312656
rect 69020 312536 69072 312588
rect 255596 312536 255648 312588
rect 370044 312536 370096 312588
rect 438860 312536 438912 312588
rect 122840 311108 122892 311160
rect 271972 311108 272024 311160
rect 400312 311108 400364 311160
rect 536840 311108 536892 311160
rect 135260 309748 135312 309800
rect 276204 309748 276256 309800
rect 406016 309748 406068 309800
rect 554780 309748 554832 309800
rect 132500 308456 132552 308508
rect 274824 308456 274876 308508
rect 74540 308388 74592 308440
rect 258356 308388 258408 308440
rect 408684 308388 408736 308440
rect 564440 308388 564492 308440
rect 207020 307096 207072 307148
rect 294604 307096 294656 307148
rect 64880 307028 64932 307080
rect 254032 307028 254084 307080
rect 381084 307028 381136 307080
rect 473360 307028 473412 307080
rect 3332 306280 3384 306332
rect 383016 306280 383068 306332
rect 379612 305668 379664 305720
rect 470600 305668 470652 305720
rect 390836 305600 390888 305652
rect 505100 305600 505152 305652
rect 209780 304308 209832 304360
rect 297456 304308 297508 304360
rect 53840 304240 53892 304292
rect 251364 304240 251416 304292
rect 413284 304240 413336 304292
rect 572812 304240 572864 304292
rect 179420 302948 179472 303000
rect 287704 302948 287756 303000
rect 15844 302880 15896 302932
rect 237656 302880 237708 302932
rect 146300 301452 146352 301504
rect 280436 301452 280488 301504
rect 393504 301452 393556 301504
rect 513380 301452 513432 301504
rect 143540 300092 143592 300144
rect 279056 300092 279108 300144
rect 397552 300092 397604 300144
rect 527180 300092 527232 300144
rect 424416 299412 424468 299464
rect 580172 299412 580224 299464
rect 361672 298732 361724 298784
rect 409880 298732 409932 298784
rect 403256 297372 403308 297424
rect 543740 297372 543792 297424
rect 402980 295944 403032 295996
rect 547880 295944 547932 295996
rect 407304 294584 407356 294636
rect 557540 294584 557592 294636
rect 2872 293904 2924 293956
rect 18604 293904 18656 293956
rect 410156 293224 410208 293276
rect 568580 293224 568632 293276
rect 154580 291796 154632 291848
rect 283196 291796 283248 291848
rect 408592 291796 408644 291848
rect 563060 291796 563112 291848
rect 136640 290436 136692 290488
rect 277584 290436 277636 290488
rect 410064 290436 410116 290488
rect 565820 290436 565872 290488
rect 157340 289144 157392 289196
rect 283104 289144 283156 289196
rect 81440 289076 81492 289128
rect 259736 289076 259788 289128
rect 411444 289076 411496 289128
rect 571984 289076 572036 289128
rect 139400 287648 139452 287700
rect 276664 287648 276716 287700
rect 397460 287648 397512 287700
rect 528560 287648 528612 287700
rect 178040 286356 178092 286408
rect 289176 286356 289228 286408
rect 354956 286356 355008 286408
rect 387800 286356 387852 286408
rect 6276 286288 6328 286340
rect 236092 286288 236144 286340
rect 376944 286288 376996 286340
rect 462320 286288 462372 286340
rect 182180 284996 182232 285048
rect 286324 284996 286376 285048
rect 356336 284996 356388 285048
rect 394700 284996 394752 285048
rect 40040 284928 40092 284980
rect 246304 284928 246356 284980
rect 285680 284928 285732 284980
rect 323216 284928 323268 284980
rect 378416 284928 378468 284980
rect 465172 284928 465224 284980
rect 184940 283636 184992 283688
rect 291384 283636 291436 283688
rect 360476 283636 360528 283688
rect 408592 283636 408644 283688
rect 35900 283568 35952 283620
rect 244924 283568 244976 283620
rect 390744 283568 390796 283620
rect 506480 283568 506532 283620
rect 195980 282208 196032 282260
rect 295524 282208 295576 282260
rect 363236 282208 363288 282260
rect 415400 282208 415452 282260
rect 20720 282140 20772 282192
rect 241796 282140 241848 282192
rect 394884 282140 394936 282192
rect 520280 282140 520332 282192
rect 200120 280848 200172 280900
rect 295984 280848 296036 280900
rect 365904 280848 365956 280900
rect 423772 280848 423824 280900
rect 121460 280780 121512 280832
rect 271144 280780 271196 280832
rect 404544 280780 404596 280832
rect 552020 280780 552072 280832
rect 296720 279624 296772 279676
rect 320824 279624 320876 279676
rect 202880 279488 202932 279540
rect 296996 279488 297048 279540
rect 365812 279488 365864 279540
rect 426440 279488 426492 279540
rect 96620 279420 96672 279472
rect 264244 279420 264296 279472
rect 405924 279420 405976 279472
rect 556160 279420 556212 279472
rect 213920 278060 213972 278112
rect 300952 278060 301004 278112
rect 372804 278060 372856 278112
rect 448520 278060 448572 278112
rect 89720 277992 89772 278044
rect 262496 277992 262548 278044
rect 412824 277992 412876 278044
rect 576124 277992 576176 278044
rect 220820 276700 220872 276752
rect 302424 276700 302476 276752
rect 85580 276632 85632 276684
rect 261116 276632 261168 276684
rect 374276 276632 374328 276684
rect 451280 276632 451332 276684
rect 227720 275340 227772 275392
rect 305184 275340 305236 275392
rect 4804 275272 4856 275324
rect 234712 275272 234764 275324
rect 375564 275272 375616 275324
rect 455420 275272 455472 275324
rect 274824 274048 274876 274100
rect 319076 274048 319128 274100
rect 129740 273912 129792 273964
rect 274640 273912 274692 273964
rect 376852 273912 376904 273964
rect 458180 273912 458232 273964
rect 431224 273164 431276 273216
rect 580172 273164 580224 273216
rect 150440 272484 150492 272536
rect 280344 272484 280396 272536
rect 359096 272484 359148 272536
rect 402980 272484 403032 272536
rect 153200 271124 153252 271176
rect 281724 271124 281776 271176
rect 381544 271124 381596 271176
rect 469220 271124 469272 271176
rect 161480 269764 161532 269816
rect 284484 269764 284536 269816
rect 383844 269764 383896 269816
rect 481640 269764 481692 269816
rect 165620 268336 165672 268388
rect 285864 268336 285916 268388
rect 383752 268336 383804 268388
rect 484400 268336 484452 268388
rect 3240 267656 3292 267708
rect 231216 267656 231268 267708
rect 222200 266976 222252 267028
rect 303712 266976 303764 267028
rect 385224 266976 385276 267028
rect 488540 266976 488592 267028
rect 168472 265616 168524 265668
rect 287244 265616 287296 265668
rect 386420 265616 386472 265668
rect 491300 265616 491352 265668
rect 172520 264188 172572 264240
rect 287152 264188 287204 264240
rect 387984 264188 388036 264240
rect 495440 264188 495492 264240
rect 183560 262828 183612 262880
rect 291292 262828 291344 262880
rect 389180 262828 389232 262880
rect 498292 262828 498344 262880
rect 292580 261536 292632 261588
rect 324596 261536 324648 261588
rect 186320 261468 186372 261520
rect 292764 261468 292816 261520
rect 354864 261468 354916 261520
rect 389180 261468 389232 261520
rect 389364 261468 389416 261520
rect 502340 261468 502392 261520
rect 190460 260108 190512 260160
rect 292856 260108 292908 260160
rect 356244 260108 356296 260160
rect 391940 260108 391992 260160
rect 392124 260108 392176 260160
rect 509240 260108 509292 260160
rect 443644 259360 443696 259412
rect 580172 259360 580224 259412
rect 193312 258748 193364 258800
rect 294144 258748 294196 258800
rect 24124 258680 24176 258732
rect 238944 258680 238996 258732
rect 364524 258680 364576 258732
rect 420920 258680 420972 258732
rect 204260 257388 204312 257440
rect 298192 257388 298244 257440
rect 22100 257320 22152 257372
rect 241704 257320 241756 257372
rect 393412 257320 393464 257372
rect 516140 257320 516192 257372
rect 208400 256028 208452 256080
rect 298376 256028 298428 256080
rect 17960 255960 18012 256012
rect 240324 255960 240376 256012
rect 357624 255960 357676 256012
rect 397460 255960 397512 256012
rect 400864 255960 400916 256012
rect 531320 255960 531372 256012
rect 3332 255212 3384 255264
rect 31024 255212 31076 255264
rect 299480 254736 299532 254788
rect 327356 254736 327408 254788
rect 211160 254600 211212 254652
rect 299756 254600 299808 254652
rect 34520 254532 34572 254584
rect 245844 254532 245896 254584
rect 357532 254532 357584 254584
rect 398932 254532 398984 254584
rect 399024 254532 399076 254584
rect 534080 254532 534132 254584
rect 303620 253376 303672 253428
rect 328736 253376 328788 253428
rect 226432 253240 226484 253292
rect 303896 253240 303948 253292
rect 33140 253172 33192 253224
rect 244464 253172 244516 253224
rect 359004 253172 359056 253224
rect 400312 253172 400364 253224
rect 400404 253172 400456 253224
rect 538220 253172 538272 253224
rect 229100 251880 229152 251932
rect 305092 251880 305144 251932
rect 29000 251812 29052 251864
rect 243084 251812 243136 251864
rect 403164 251812 403216 251864
rect 545120 251812 545172 251864
rect 276204 250588 276256 250640
rect 318984 250588 319036 250640
rect 133880 250452 133932 250504
rect 276112 250452 276164 250504
rect 404452 250452 404504 250504
rect 547972 250452 548024 250504
rect 233240 249092 233292 249144
rect 306472 249092 306524 249144
rect 16580 249024 16632 249076
rect 233976 249024 234028 249076
rect 409972 249024 410024 249076
rect 569960 249024 570012 249076
rect 140780 247664 140832 247716
rect 277492 247664 277544 247716
rect 367284 247664 367336 247716
rect 432052 247664 432104 247716
rect 143632 246304 143684 246356
rect 278964 246304 279016 246356
rect 385132 246304 385184 246356
rect 485780 246304 485832 246356
rect 422944 245556 422996 245608
rect 580172 245556 580224 245608
rect 147680 244876 147732 244928
rect 280252 244876 280304 244928
rect 386512 243584 386564 243636
rect 151820 243516 151872 243568
rect 281632 243516 281684 243568
rect 353484 243516 353536 243568
rect 386420 243516 386472 243568
rect 492680 243516 492732 243568
rect 158720 242156 158772 242208
rect 283012 242156 283064 242208
rect 387892 242156 387944 242208
rect 496820 242156 496872 242208
rect 3240 241408 3292 241460
rect 232596 241408 232648 241460
rect 389272 240728 389324 240780
rect 499580 240728 499632 240780
rect 167000 239368 167052 239420
rect 285772 239368 285824 239420
rect 390652 239368 390704 239420
rect 503720 239368 503772 239420
rect 180800 238008 180852 238060
rect 290004 238008 290056 238060
rect 392032 238008 392084 238060
rect 510620 238008 510672 238060
rect 187700 236648 187752 236700
rect 292672 236648 292724 236700
rect 394792 236648 394844 236700
rect 517520 236648 517572 236700
rect 191840 235220 191892 235272
rect 294052 235220 294104 235272
rect 396264 235220 396316 235272
rect 521660 235220 521712 235272
rect 131120 233860 131172 233912
rect 274732 233860 274784 233912
rect 396172 233860 396224 233912
rect 524420 233860 524472 233912
rect 438124 233180 438176 233232
rect 579620 233180 579672 233232
rect 201592 232500 201644 232552
rect 296812 232500 296864 232552
rect 209872 231072 209924 231124
rect 299664 231072 299716 231124
rect 401784 231072 401836 231124
rect 539600 231072 539652 231124
rect 212540 229712 212592 229764
rect 299572 229712 299624 229764
rect 401692 229712 401744 229764
rect 542360 229712 542412 229764
rect 142160 228352 142212 228404
rect 278872 228352 278924 228404
rect 403072 228352 403124 228404
rect 546500 228352 546552 228404
rect 100760 226992 100812 227044
rect 265164 226992 265216 227044
rect 405832 226992 405884 227044
rect 553400 226992 553452 227044
rect 103520 225564 103572 225616
rect 266544 225564 266596 225616
rect 407212 225564 407264 225616
rect 560300 225564 560352 225616
rect 44180 224204 44232 224256
rect 248604 224204 248656 224256
rect 411352 224204 411404 224256
rect 574100 224204 574152 224256
rect 13084 222844 13136 222896
rect 237564 222844 237616 222896
rect 48320 221416 48372 221468
rect 249984 221416 250036 221468
rect 52460 220056 52512 220108
rect 249892 220056 249944 220108
rect 442264 219376 442316 219428
rect 580172 219376 580224 219428
rect 59360 218696 59412 218748
rect 252744 218696 252796 218748
rect 62120 217268 62172 217320
rect 251824 217268 251876 217320
rect 66260 215908 66312 215960
rect 255504 215908 255556 215960
rect 2780 214956 2832 215008
rect 4896 214956 4948 215008
rect 84200 214548 84252 214600
rect 261024 214548 261076 214600
rect 86960 213188 87012 213240
rect 260932 213188 260984 213240
rect 98000 211760 98052 211812
rect 265072 211760 265124 211812
rect 104900 210400 104952 210452
rect 266452 210400 266504 210452
rect 30380 209040 30432 209092
rect 244372 209040 244424 209092
rect 41420 207612 41472 207664
rect 247224 207612 247276 207664
rect 421564 206932 421616 206984
rect 580172 206932 580224 206984
rect 56600 206252 56652 206304
rect 252652 206252 252704 206304
rect 63500 204892 63552 204944
rect 254216 204892 254268 204944
rect 67640 203532 67692 203584
rect 255412 203532 255464 203584
rect 3332 202784 3384 202836
rect 11796 202784 11848 202836
rect 70400 202104 70452 202156
rect 256884 202104 256936 202156
rect 77300 200744 77352 200796
rect 258264 200744 258316 200796
rect 88340 199384 88392 199436
rect 262404 199384 262456 199436
rect 92480 197956 92532 198008
rect 262312 197956 262364 198008
rect 95240 196596 95292 196648
rect 263784 196596 263836 196648
rect 106280 195236 106332 195288
rect 267924 195236 267976 195288
rect 429844 193128 429896 193180
rect 580172 193128 580224 193180
rect 3148 188980 3200 189032
rect 40684 188980 40736 189032
rect 440884 179324 440936 179376
rect 580172 179324 580224 179376
rect 420184 166948 420236 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 229744 164160 229796 164212
rect 428464 153144 428516 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 13176 150356 13228 150408
rect 439504 139340 439556 139392
rect 580172 139340 580224 139392
rect 435364 126896 435416 126948
rect 579620 126896 579672 126948
rect 427084 113092 427136 113144
rect 580172 113092 580224 113144
rect 7656 111052 7708 111104
rect 234804 111052 234856 111104
rect 3240 110984 3292 111036
rect 7564 110984 7616 111036
rect 436744 100648 436796 100700
rect 579712 100648 579764 100700
rect 3240 97928 3292 97980
rect 14464 97928 14516 97980
rect 14556 97248 14608 97300
rect 237472 97248 237524 97300
rect 418804 86912 418856 86964
rect 579988 86912 580040 86964
rect 3332 85484 3384 85536
rect 21364 85484 21416 85536
rect 425704 73108 425756 73160
rect 580172 73108 580224 73160
rect 3332 71680 3384 71732
rect 233884 71680 233936 71732
rect 27620 68280 27672 68332
rect 242992 68280 243044 68332
rect 44272 64132 44324 64184
rect 248512 64132 248564 64184
rect 99380 62772 99432 62824
rect 265256 62772 265308 62824
rect 52552 61344 52604 61396
rect 251272 61344 251324 61396
rect 432604 60664 432656 60716
rect 579804 60664 579856 60716
rect 102232 59984 102284 60036
rect 266636 59984 266688 60036
rect 3332 59304 3384 59356
rect 28264 59304 28316 59356
rect 160192 58624 160244 58676
rect 284392 58624 284444 58676
rect 155960 57196 156012 57248
rect 282920 57196 282972 57248
rect 151912 55836 151964 55888
rect 281540 55836 281592 55888
rect 135352 54476 135404 54528
rect 276020 54476 276072 54528
rect 149060 53048 149112 53100
rect 280160 53048 280212 53100
rect 69112 51688 69164 51740
rect 255320 51688 255372 51740
rect 255412 51688 255464 51740
rect 313372 51688 313424 51740
rect 396080 51688 396132 51740
rect 523040 51688 523092 51740
rect 49700 50328 49752 50380
rect 249800 50328 249852 50380
rect 251272 50328 251324 50380
rect 312084 50328 312136 50380
rect 244372 48968 244424 49020
rect 310704 48968 310756 49020
rect 237472 47540 237524 47592
rect 307852 47540 307904 47592
rect 417424 46860 417476 46912
rect 580172 46860 580224 46912
rect 234620 46180 234672 46232
rect 305644 46180 305696 46232
rect 363144 46180 363196 46232
rect 416780 46180 416832 46232
rect 230480 44820 230532 44872
rect 305000 44820 305052 44872
rect 216680 43392 216732 43444
rect 300860 43392 300912 43444
rect 198740 42032 198792 42084
rect 295432 42032 295484 42084
rect 194600 40672 194652 40724
rect 294236 40672 294288 40724
rect 185032 39312 185084 39364
rect 291476 39312 291528 39364
rect 310704 39312 310756 39364
rect 330116 39312 330168 39364
rect 169760 37884 169812 37936
rect 287336 37884 287388 37936
rect 138020 36524 138072 36576
rect 277676 36524 277728 36576
rect 282920 36524 282972 36576
rect 321836 36524 321888 36576
rect 85672 35164 85724 35216
rect 260840 35164 260892 35216
rect 267924 35164 267976 35216
rect 317604 35164 317656 35216
rect 73160 33736 73212 33788
rect 256792 33736 256844 33788
rect 258264 33736 258316 33788
rect 314752 33736 314804 33788
rect 2780 32444 2832 32496
rect 6184 32444 6236 32496
rect 55220 32376 55272 32428
rect 251180 32376 251232 32428
rect 251364 32376 251416 32428
rect 311992 32376 312044 32428
rect 358912 32376 358964 32428
rect 404452 32376 404504 32428
rect 411260 32376 411312 32428
rect 571340 32376 571392 32428
rect 247224 31016 247276 31068
rect 310612 31016 310664 31068
rect 356152 31016 356204 31068
rect 393412 31016 393464 31068
rect 242992 29588 243044 29640
rect 309324 29588 309376 29640
rect 354772 29588 354824 29640
rect 390744 29588 390796 29640
rect 400220 29588 400272 29640
rect 535460 29588 535512 29640
rect 240324 28228 240376 28280
rect 309232 28228 309284 28280
rect 350632 28228 350684 28280
rect 375564 28228 375616 28280
rect 393320 28228 393372 28280
rect 514852 28228 514904 28280
rect 262312 26936 262364 26988
rect 316224 26936 316276 26988
rect 218060 26868 218112 26920
rect 298744 26868 298796 26920
rect 347964 26868 348016 26920
rect 365812 26868 365864 26920
rect 390560 26868 390612 26920
rect 506572 26868 506624 26920
rect 162860 25576 162912 25628
rect 284576 25576 284628 25628
rect 284392 25508 284444 25560
rect 323124 25508 323176 25560
rect 360384 25508 360436 25560
rect 407212 25508 407264 25560
rect 408500 25508 408552 25560
rect 564532 25508 564584 25560
rect 353392 24216 353444 24268
rect 385132 24216 385184 24268
rect 259736 24148 259788 24200
rect 307116 24148 307168 24200
rect 126980 24080 127032 24132
rect 273352 24080 273404 24132
rect 281540 24080 281592 24132
rect 321744 24080 321796 24132
rect 385040 24080 385092 24132
rect 490012 24080 490064 24132
rect 248512 22788 248564 22840
rect 310796 22788 310848 22840
rect 60832 22720 60884 22772
rect 252836 22720 252888 22772
rect 263784 22720 263836 22772
rect 316132 22720 316184 22772
rect 356060 22720 356112 22772
rect 396080 22720 396132 22772
rect 398840 22720 398892 22772
rect 531412 22720 531464 22772
rect 256792 21428 256844 21480
rect 313464 21428 313516 21480
rect 144920 21360 144972 21412
rect 278780 21360 278832 21412
rect 352104 21360 352156 21412
rect 382464 21360 382516 21412
rect 383660 21360 383712 21412
rect 481732 21360 481784 21412
rect 3516 20612 3568 20664
rect 414940 20612 414992 20664
rect 360292 18708 360344 18760
rect 405832 18708 405884 18760
rect 289820 18640 289872 18692
rect 315304 18640 315356 18692
rect 37280 18572 37332 18624
rect 245752 18572 245804 18624
rect 249800 18572 249852 18624
rect 297364 18572 297416 18624
rect 405740 18572 405792 18624
rect 556252 18572 556304 18624
rect 243084 17280 243136 17332
rect 302976 17280 303028 17332
rect 358084 17280 358136 17332
rect 372804 17280 372856 17332
rect 241704 17212 241756 17264
rect 309416 17212 309468 17264
rect 346584 17212 346636 17264
rect 360292 17212 360344 17264
rect 370504 17212 370556 17264
rect 412824 17212 412876 17264
rect 260656 15920 260708 15972
rect 291844 15920 291896 15972
rect 116400 15852 116452 15904
rect 270684 15852 270736 15904
rect 279056 15852 279108 15904
rect 319444 15852 319496 15904
rect 358820 15852 358872 15904
rect 402520 15852 402572 15904
rect 404360 15852 404412 15904
rect 550272 15852 550324 15904
rect 112352 14764 112404 14816
rect 269304 14764 269356 14816
rect 109040 14696 109092 14748
rect 267832 14696 267884 14748
rect 93860 14628 93912 14680
rect 263692 14628 263744 14680
rect 91560 14560 91612 14612
rect 262220 14560 262272 14612
rect 80888 14492 80940 14544
rect 259644 14492 259696 14544
rect 77392 14424 77444 14476
rect 258172 14424 258224 14476
rect 267740 14424 267792 14476
rect 313924 14424 313976 14476
rect 352012 14424 352064 14476
rect 381176 14424 381228 14476
rect 407120 14424 407172 14476
rect 559288 14424 559340 14476
rect 313832 13948 313884 14000
rect 318064 13948 318116 14000
rect 118792 13336 118844 13388
rect 270592 13336 270644 13388
rect 114744 13268 114796 13320
rect 270776 13268 270828 13320
rect 111616 13200 111668 13252
rect 269212 13200 269264 13252
rect 108120 13132 108172 13184
rect 268108 13132 268160 13184
rect 350540 13132 350592 13184
rect 377312 13132 377364 13184
rect 93952 13064 94004 13116
rect 263600 13064 263652 13116
rect 270776 13064 270828 13116
rect 317512 13064 317564 13116
rect 363052 13064 363104 13116
rect 415492 13064 415544 13116
rect 417516 13064 417568 13116
rect 541992 13064 542044 13116
rect 160100 11772 160152 11824
rect 161296 11772 161348 11824
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 226340 11772 226392 11824
rect 227536 11772 227588 11824
rect 254216 11772 254268 11824
rect 307024 11772 307076 11824
rect 349344 11772 349396 11824
rect 374276 11772 374328 11824
rect 12992 11704 13044 11756
rect 238852 11704 238904 11756
rect 239312 11704 239364 11756
rect 301504 11704 301556 11756
rect 307944 11704 307996 11756
rect 330024 11704 330076 11756
rect 373264 11704 373316 11756
rect 414020 11704 414072 11756
rect 424324 11704 424376 11756
rect 523132 11704 523184 11756
rect 372620 10820 372672 10872
rect 445760 10820 445812 10872
rect 372712 10752 372764 10804
rect 448612 10752 448664 10804
rect 374184 10684 374236 10736
rect 453304 10684 453356 10736
rect 375472 10616 375524 10668
rect 456892 10616 456944 10668
rect 376760 10548 376812 10600
rect 459928 10548 459980 10600
rect 378324 10480 378376 10532
rect 463976 10480 464028 10532
rect 173900 10412 173952 10464
rect 288532 10412 288584 10464
rect 378232 10412 378284 10464
rect 467472 10412 467524 10464
rect 83280 10344 83332 10396
rect 259552 10344 259604 10396
rect 288992 10344 289044 10396
rect 323032 10344 323084 10396
rect 345112 10344 345164 10396
rect 357532 10344 357584 10396
rect 380992 10344 381044 10396
rect 474096 10344 474148 10396
rect 79232 10276 79284 10328
rect 259460 10276 259512 10328
rect 264980 10276 265032 10328
rect 302884 10276 302936 10328
rect 349252 10276 349304 10328
rect 371516 10276 371568 10328
rect 382372 10276 382424 10328
rect 478144 10276 478196 10328
rect 209688 9596 209740 9648
rect 210976 9596 211028 9648
rect 253480 9052 253532 9104
rect 312176 9052 312228 9104
rect 76196 8984 76248 9036
rect 258080 8984 258132 9036
rect 349160 8984 349212 9036
rect 370596 8984 370648 9036
rect 72608 8916 72660 8968
rect 256700 8916 256752 8968
rect 261760 8916 261812 8968
rect 314844 8916 314896 8968
rect 317328 8916 317380 8968
rect 332784 8916 332836 8968
rect 351920 8916 351972 8968
rect 379980 8916 380032 8968
rect 387064 8916 387116 8968
rect 398840 8916 398892 8968
rect 412732 8916 412784 8968
rect 577412 8916 577464 8968
rect 377404 8236 377456 8288
rect 378876 8236 378928 8288
rect 272432 7692 272484 7744
rect 318892 7692 318944 7744
rect 197912 7624 197964 7676
rect 295340 7624 295392 7676
rect 347872 7624 347924 7676
rect 367008 7624 367060 7676
rect 176752 7556 176804 7608
rect 288716 7556 288768 7608
rect 310244 7556 310296 7608
rect 329932 7556 329984 7608
rect 347780 7556 347832 7608
rect 369400 7556 369452 7608
rect 380900 7556 380952 7608
rect 476948 7556 477000 7608
rect 3516 6468 3568 6520
rect 8944 6468 8996 6520
rect 367192 6468 367244 6520
rect 430856 6468 430908 6520
rect 368664 6400 368716 6452
rect 434444 6400 434496 6452
rect 369952 6332 370004 6384
rect 437940 6332 437992 6384
rect 235816 6264 235868 6316
rect 306564 6264 306616 6316
rect 371332 6264 371384 6316
rect 441528 6264 441580 6316
rect 237012 6196 237064 6248
rect 304264 6196 304316 6248
rect 345020 6196 345072 6248
rect 359924 6196 359976 6248
rect 371424 6196 371476 6248
rect 445024 6196 445076 6248
rect 128176 6128 128228 6180
rect 231124 6128 231176 6180
rect 306748 6128 306800 6180
rect 328644 6128 328696 6180
rect 346492 6128 346544 6180
rect 364616 6128 364668 6180
rect 412640 6128 412692 6180
rect 576308 6128 576360 6180
rect 366364 5516 366416 5568
rect 368204 5516 368256 5568
rect 303160 5040 303212 5092
rect 328552 5040 328604 5092
rect 299664 4972 299716 5024
rect 327264 4972 327316 5024
rect 296076 4904 296128 4956
rect 325792 4904 325844 4956
rect 351184 4904 351236 4956
rect 356336 4904 356388 4956
rect 278320 4836 278372 4888
rect 320364 4836 320416 4888
rect 353300 4836 353352 4888
rect 383568 4836 383620 4888
rect 218152 4768 218204 4820
rect 228364 4768 228416 4820
rect 246396 4768 246448 4820
rect 289084 4768 289136 4820
rect 292580 4768 292632 4820
rect 324504 4768 324556 4820
rect 354680 4768 354732 4820
rect 391848 4768 391900 4820
rect 401600 4768 401652 4820
rect 540796 4768 540848 4820
rect 382924 4496 382976 4548
rect 384764 4496 384816 4548
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 176660 4156 176712 4208
rect 177856 4156 177908 4208
rect 345664 4156 345716 4208
rect 352840 4156 352892 4208
rect 46664 4088 46716 4140
rect 248696 4088 248748 4140
rect 305552 4088 305604 4140
rect 328460 4088 328512 4140
rect 332692 4088 332744 4140
rect 336924 4088 336976 4140
rect 341156 4088 341208 4140
rect 345756 4088 345808 4140
rect 367100 4088 367152 4140
rect 429660 4088 429712 4140
rect 43076 4020 43128 4072
rect 247316 4020 247368 4072
rect 301964 4020 302016 4072
rect 327080 4020 327132 4072
rect 39580 3952 39632 4004
rect 247132 3952 247184 4004
rect 298468 3952 298520 4004
rect 327172 3952 327224 4004
rect 2872 3884 2924 3936
rect 7656 3884 7708 3936
rect 35992 3884 36044 3936
rect 245936 3884 245988 3936
rect 294880 3884 294932 3936
rect 325884 3884 325936 3936
rect 326804 3884 326856 3936
rect 335544 4020 335596 4072
rect 340972 4020 341024 4072
rect 346952 4020 347004 4072
rect 368572 4020 368624 4072
rect 433248 4020 433300 4072
rect 333888 3952 333940 4004
rect 337108 3952 337160 4004
rect 368480 3952 368532 4004
rect 436744 3952 436796 4004
rect 328000 3884 328052 3936
rect 335360 3884 335412 3936
rect 342536 3884 342588 3936
rect 348056 3884 348108 3936
rect 369860 3884 369912 3936
rect 440332 3884 440384 3936
rect 32404 3816 32456 3868
rect 244280 3816 244332 3868
rect 291384 3816 291436 3868
rect 324412 3816 324464 3868
rect 329196 3816 329248 3868
rect 335636 3816 335688 3868
rect 342628 3816 342680 3868
rect 350448 3816 350500 3868
rect 371240 3816 371292 3868
rect 443828 3816 443880 3868
rect 28908 3748 28960 3800
rect 242900 3748 242952 3800
rect 287796 3748 287848 3800
rect 322940 3748 322992 3800
rect 325608 3748 325660 3800
rect 335452 3748 335504 3800
rect 374184 3748 374236 3800
rect 450912 3748 450964 3800
rect 576124 3748 576176 3800
rect 578608 3748 578660 3800
rect 14740 3680 14792 3732
rect 24124 3680 24176 3732
rect 25320 3680 25372 3732
rect 241520 3680 241572 3732
rect 284300 3680 284352 3732
rect 321560 3680 321612 3732
rect 323308 3680 323360 3732
rect 334164 3680 334216 3732
rect 342444 3680 342496 3732
rect 349252 3680 349304 3732
rect 375380 3680 375432 3732
rect 458088 3680 458140 3732
rect 8760 3612 8812 3664
rect 13084 3612 13136 3664
rect 24216 3612 24268 3664
rect 241612 3612 241664 3664
rect 280712 3612 280764 3664
rect 321652 3612 321704 3664
rect 322112 3612 322164 3664
rect 334072 3612 334124 3664
rect 346400 3612 346452 3664
rect 362316 3612 362368 3664
rect 378140 3612 378192 3664
rect 465172 3612 465224 3664
rect 6460 3544 6512 3596
rect 10324 3544 10376 3596
rect 19432 3544 19484 3596
rect 240232 3544 240284 3596
rect 242900 3544 242952 3596
rect 243084 3544 243136 3596
rect 251272 3544 251324 3596
rect 252376 3544 252428 3596
rect 273628 3544 273680 3596
rect 318800 3544 318852 3596
rect 319720 3544 319772 3596
rect 332600 3544 332652 3596
rect 342352 3544 342404 3596
rect 351644 3544 351696 3596
rect 360200 3544 360252 3596
rect 408408 3544 408460 3596
rect 414204 3544 414256 3596
rect 582196 3544 582248 3596
rect 572 3476 624 3528
rect 3424 3476 3476 3528
rect 12348 3476 12400 3528
rect 15844 3476 15896 3528
rect 20628 3476 20680 3528
rect 240416 3476 240468 3528
rect 266544 3476 266596 3528
rect 316316 3476 316368 3528
rect 318524 3476 318576 3528
rect 332508 3476 332560 3528
rect 337476 3476 337528 3528
rect 338396 3476 338448 3528
rect 338672 3476 338724 3528
rect 339592 3476 339644 3528
rect 339684 3476 339736 3528
rect 340972 3476 341024 3528
rect 343732 3476 343784 3528
rect 354036 3476 354088 3528
rect 357440 3476 357492 3528
rect 358728 3476 358780 3528
rect 374000 3476 374052 3528
rect 375288 3476 375340 3528
rect 379520 3476 379572 3528
rect 472256 3476 472308 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 1676 3408 1728 3460
rect 4804 3408 4856 3460
rect 9956 3408 10008 3460
rect 14556 3408 14608 3460
rect 15936 3408 15988 3460
rect 238760 3408 238812 3460
rect 299480 3408 299532 3460
rect 300768 3408 300820 3460
rect 316224 3408 316276 3460
rect 331496 3408 331548 3460
rect 343640 3408 343692 3460
rect 355232 3408 355284 3460
rect 361580 3408 361632 3460
rect 411904 3408 411956 3460
rect 415400 3408 415452 3460
rect 416688 3408 416740 3460
rect 416780 3408 416832 3460
rect 581000 3408 581052 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 77300 3340 77352 3392
rect 78220 3340 78272 3392
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 7656 3272 7708 3324
rect 11704 3272 11756 3324
rect 114008 3272 114060 3324
rect 269120 3340 269172 3392
rect 309048 3340 309100 3392
rect 329840 3340 329892 3392
rect 341064 3340 341116 3392
rect 344560 3340 344612 3392
rect 365720 3340 365772 3392
rect 426164 3340 426216 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 121092 3272 121144 3324
rect 272156 3272 272208 3324
rect 312636 3272 312688 3324
rect 331312 3272 331364 3324
rect 364432 3272 364484 3324
rect 422576 3272 422628 3324
rect 124680 3204 124732 3256
rect 273444 3204 273496 3256
rect 315028 3204 315080 3256
rect 331404 3204 331456 3256
rect 218060 3136 218112 3188
rect 219256 3136 219308 3188
rect 270040 3136 270092 3188
rect 317696 3136 317748 3188
rect 330392 3136 330444 3188
rect 336832 3204 336884 3256
rect 364340 3204 364392 3256
rect 418988 3204 419040 3256
rect 336280 3136 336332 3188
rect 338212 3136 338264 3188
rect 398932 3136 398984 3188
rect 400128 3136 400180 3188
rect 414112 3136 414164 3188
rect 416780 3136 416832 3188
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 4068 2864 4120 2916
rect 6276 2864 6328 2916
rect 423680 960 423732 1012
rect 424968 960 425020 1012
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3344 618322 3372 619103
rect 3332 618316 3384 618322
rect 3332 618258 3384 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3436 460193 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3528 465746 3556 632023
rect 3606 580000 3662 580009
rect 3606 579935 3662 579944
rect 3620 465882 3648 579935
rect 3698 527912 3754 527921
rect 3698 527847 3754 527856
rect 3712 466018 3740 527847
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3712 465990 3832 466018
rect 3620 465854 3740 465882
rect 3528 465718 3648 465746
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3620 460426 3648 465718
rect 3608 460420 3660 460426
rect 3608 460362 3660 460368
rect 3712 460358 3740 465854
rect 3700 460352 3752 460358
rect 3700 460294 3752 460300
rect 3804 460290 3832 465990
rect 3792 460284 3844 460290
rect 3792 460226 3844 460232
rect 3896 460222 3924 475623
rect 4896 460964 4948 460970
rect 4896 460906 4948 460912
rect 3884 460216 3936 460222
rect 3422 460184 3478 460193
rect 3884 460158 3936 460164
rect 3422 460119 3478 460128
rect 3424 458856 3476 458862
rect 3424 458798 3476 458804
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3436 358465 3464 458798
rect 3608 458244 3660 458250
rect 3608 458186 3660 458192
rect 3516 457496 3568 457502
rect 3516 457438 3568 457444
rect 3528 397497 3556 457438
rect 3620 423609 3648 458186
rect 3606 423600 3662 423609
rect 3606 423535 3662 423544
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3516 372564 3568 372570
rect 3516 372506 3568 372512
rect 3528 371385 3556 372506
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3424 334620 3476 334626
rect 3424 334562 3476 334568
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2872 293956 2924 293962
rect 2872 293898 2924 293904
rect 2884 293185 2912 293898
rect 2870 293176 2926 293185
rect 2870 293111 2926 293120
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3332 255264 3384 255270
rect 3332 255206 3384 255212
rect 3344 254153 3372 255206
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 2780 215008 2832 215014
rect 2778 214976 2780 214985
rect 2832 214976 2834 214985
rect 2778 214911 2834 214920
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3240 111036 3292 111042
rect 3240 110978 3292 110984
rect 3252 110673 3280 110978
rect 3238 110664 3294 110673
rect 3238 110599 3294 110608
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3332 59356 3384 59362
rect 3332 59298 3384 59304
rect 3344 58585 3372 59298
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 2780 32496 2832 32502
rect 2778 32464 2780 32473
rect 2832 32464 2834 32473
rect 2778 32399 2834 32408
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3878
rect 3436 3534 3464 334562
rect 3516 320136 3568 320142
rect 3516 320078 3568 320084
rect 3528 319297 3556 320078
rect 3514 319288 3570 319297
rect 3514 319223 3570 319232
rect 3606 316704 3662 316713
rect 3606 316639 3662 316648
rect 3514 313984 3570 313993
rect 3514 313919 3570 313928
rect 3528 45529 3556 313919
rect 3620 136785 3648 316639
rect 4804 275324 4856 275330
rect 4804 275266 4856 275272
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3516 6520 3568 6526
rect 3514 6488 3516 6497
rect 3568 6488 3570 6497
rect 3514 6423 3570 6432
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 4816 3466 4844 275266
rect 4908 215014 4936 460906
rect 40052 460329 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 104912 460494 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 460698 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700602 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700596 154172 700602
rect 154120 700538 154172 700544
rect 169772 468518 169800 702406
rect 169760 468512 169812 468518
rect 169760 468454 169812 468460
rect 201512 460834 201540 702986
rect 218992 700738 219020 703520
rect 218980 700732 219032 700738
rect 218980 700674 219032 700680
rect 235184 698970 235212 703520
rect 235172 698964 235224 698970
rect 235172 698906 235224 698912
rect 267660 697610 267688 703520
rect 283852 700874 283880 703520
rect 283840 700868 283892 700874
rect 283840 700810 283892 700816
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 226984 462528 227036 462534
rect 226984 462470 227036 462476
rect 201500 460828 201552 460834
rect 201500 460770 201552 460776
rect 136640 460692 136692 460698
rect 136640 460634 136692 460640
rect 104900 460488 104952 460494
rect 104900 460430 104952 460436
rect 40038 460320 40094 460329
rect 40038 460255 40094 460264
rect 226996 411262 227024 462470
rect 233976 461372 234028 461378
rect 233976 461314 234028 461320
rect 228364 461100 228416 461106
rect 228364 461042 228416 461048
rect 226984 411256 227036 411262
rect 226984 411198 227036 411204
rect 228376 346390 228404 461042
rect 229744 461032 229796 461038
rect 229744 460974 229796 460980
rect 228364 346384 228416 346390
rect 228364 346326 228416 346332
rect 7562 337376 7618 337385
rect 7562 337311 7618 337320
rect 6182 333296 6238 333305
rect 6182 333231 6238 333240
rect 4896 215008 4948 215014
rect 4896 214950 4948 214956
rect 6196 32502 6224 333231
rect 6276 286340 6328 286346
rect 6276 286282 6328 286288
rect 6184 32496 6236 32502
rect 6184 32438 6236 32444
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4080 480 4108 2858
rect 5276 480 5304 3295
rect 6288 2922 6316 286282
rect 7576 111042 7604 337311
rect 228364 336320 228416 336326
rect 228364 336262 228416 336268
rect 117320 336252 117372 336258
rect 117320 336194 117372 336200
rect 110420 336184 110472 336190
rect 110420 336126 110472 336132
rect 102140 336116 102192 336122
rect 102140 336058 102192 336064
rect 10324 336048 10376 336054
rect 10324 335990 10376 335996
rect 8942 311128 8998 311137
rect 8942 311063 8998 311072
rect 7656 111104 7708 111110
rect 7656 111046 7708 111052
rect 7564 111036 7616 111042
rect 7564 110978 7616 110984
rect 7668 3942 7696 111046
rect 8956 6526 8984 311063
rect 8944 6520 8996 6526
rect 8944 6462 8996 6468
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6472 480 6500 3538
rect 7656 3324 7708 3330
rect 7656 3266 7708 3272
rect 7668 480 7696 3266
rect 8772 480 8800 3606
rect 10336 3602 10364 335990
rect 46940 331900 46992 331906
rect 46940 331842 46992 331848
rect 11704 326392 11756 326398
rect 11704 326334 11756 326340
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11150 3496 11206 3505
rect 9956 3460 10008 3466
rect 11150 3431 11206 3440
rect 9956 3402 10008 3408
rect 9968 480 9996 3402
rect 11164 480 11192 3431
rect 11716 3330 11744 326334
rect 26240 323604 26292 323610
rect 26240 323546 26292 323552
rect 18602 320784 18658 320793
rect 18602 320719 18658 320728
rect 15844 302932 15896 302938
rect 15844 302874 15896 302880
rect 11794 297392 11850 297401
rect 11794 297327 11850 297336
rect 11808 202842 11836 297327
rect 13174 296032 13230 296041
rect 13174 295967 13230 295976
rect 13084 222896 13136 222902
rect 13084 222838 13136 222844
rect 11796 202836 11848 202842
rect 11796 202778 11848 202784
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 13004 3482 13032 11698
rect 13096 3670 13124 222838
rect 13188 150414 13216 295967
rect 14462 294536 14518 294545
rect 14462 294471 14518 294480
rect 13176 150408 13228 150414
rect 13176 150350 13228 150356
rect 14476 97986 14504 294471
rect 14464 97980 14516 97986
rect 14464 97922 14516 97928
rect 14556 97300 14608 97306
rect 14556 97242 14608 97248
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 11704 3324 11756 3330
rect 11704 3266 11756 3272
rect 12360 480 12388 3470
rect 13004 3454 13584 3482
rect 14568 3466 14596 97242
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 13556 480 13584 3454
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14752 480 14780 3674
rect 15856 3534 15884 302874
rect 18616 293962 18644 320719
rect 21362 315344 21418 315353
rect 21362 315279 21418 315288
rect 18604 293956 18656 293962
rect 18604 293898 18656 293904
rect 20720 282192 20772 282198
rect 20720 282134 20772 282140
rect 17960 256012 18012 256018
rect 17960 255954 18012 255960
rect 16580 249076 16632 249082
rect 16580 249018 16632 249024
rect 16592 16574 16620 249018
rect 16592 16546 17080 16574
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 480 15976 3402
rect 17052 480 17080 16546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 255954
rect 20732 16574 20760 282134
rect 21376 85542 21404 315279
rect 24124 258732 24176 258738
rect 24124 258674 24176 258680
rect 22100 257372 22152 257378
rect 22100 257314 22152 257320
rect 21364 85536 21416 85542
rect 21364 85478 21416 85484
rect 22112 16574 22140 257314
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19444 480 19472 3538
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 480 20668 3470
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24136 3738 24164 258674
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 480 24256 3606
rect 25332 480 25360 3674
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 323546
rect 40682 318064 40738 318073
rect 40682 317999 40738 318008
rect 31022 298752 31078 298761
rect 31022 298687 31078 298696
rect 28262 293176 28318 293185
rect 28262 293111 28318 293120
rect 27620 68332 27672 68338
rect 27620 68274 27672 68280
rect 27632 16574 27660 68274
rect 28276 59362 28304 293111
rect 31036 255270 31064 298687
rect 40040 284980 40092 284986
rect 40040 284922 40092 284928
rect 35900 283620 35952 283626
rect 35900 283562 35952 283568
rect 31024 255264 31076 255270
rect 31024 255206 31076 255212
rect 34520 254584 34572 254590
rect 34520 254526 34572 254532
rect 33140 253224 33192 253230
rect 33140 253166 33192 253172
rect 29000 251864 29052 251870
rect 29000 251806 29052 251812
rect 28264 59356 28316 59362
rect 28264 59298 28316 59304
rect 29012 16574 29040 251806
rect 30380 209092 30432 209098
rect 30380 209034 30432 209040
rect 30392 16574 30420 209034
rect 33152 16574 33180 253166
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 16546
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 32404 3868 32456 3874
rect 32404 3810 32456 3816
rect 32416 480 32444 3810
rect 33612 480 33640 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 254526
rect 35912 16574 35940 283562
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37292 16574 37320 18566
rect 40052 16574 40080 284922
rect 40696 189038 40724 317999
rect 44180 224256 44232 224262
rect 44180 224198 44232 224204
rect 41420 207664 41472 207670
rect 41420 207606 41472 207612
rect 40684 189032 40736 189038
rect 40684 188974 40736 188980
rect 41432 16574 41460 207606
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35992 3936 36044 3942
rect 35992 3878 36044 3884
rect 36004 480 36032 3878
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 39580 4004 39632 4010
rect 39580 3946 39632 3952
rect 39592 480 39620 3946
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 44192 6914 44220 224198
rect 44272 64184 44324 64190
rect 44272 64126 44324 64132
rect 44284 16574 44312 64126
rect 46952 16574 46980 331842
rect 57980 330540 58032 330546
rect 57980 330482 58032 330488
rect 51080 322244 51132 322250
rect 51080 322186 51132 322192
rect 48320 221468 48372 221474
rect 48320 221410 48372 221416
rect 48332 16574 48360 221410
rect 49700 50380 49752 50386
rect 49700 50322 49752 50328
rect 49712 16574 49740 50322
rect 44284 16546 45048 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43088 480 43116 4014
rect 44284 480 44312 6886
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46664 4140 46716 4146
rect 46664 4082 46716 4088
rect 46676 480 46704 4082
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 322186
rect 53840 304292 53892 304298
rect 53840 304234 53892 304240
rect 52460 220108 52512 220114
rect 52460 220050 52512 220056
rect 52472 6914 52500 220050
rect 52552 61396 52604 61402
rect 52552 61338 52604 61344
rect 52564 16574 52592 61338
rect 53852 16574 53880 304234
rect 56600 206304 56652 206310
rect 56600 206246 56652 206252
rect 55220 32428 55272 32434
rect 55220 32370 55272 32376
rect 55232 16574 55260 32370
rect 56612 16574 56640 206246
rect 57992 16574 58020 330482
rect 60740 329112 60792 329118
rect 60740 329054 60792 329060
rect 59360 218748 59412 218754
rect 59360 218690 59412 218696
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 218690
rect 60752 3398 60780 329054
rect 69020 312588 69072 312594
rect 69020 312530 69072 312536
rect 64880 307080 64932 307086
rect 64880 307022 64932 307028
rect 62120 217320 62172 217326
rect 62120 217262 62172 217268
rect 60832 22772 60884 22778
rect 60832 22714 60884 22720
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 22714
rect 62132 16574 62160 217262
rect 63500 204944 63552 204950
rect 63500 204886 63552 204892
rect 63512 16574 63540 204886
rect 64892 16574 64920 307022
rect 66260 215960 66312 215966
rect 66260 215902 66312 215908
rect 66272 16574 66300 215902
rect 67640 203584 67692 203590
rect 67640 203526 67692 203532
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 203526
rect 69032 6914 69060 312530
rect 74540 308440 74592 308446
rect 74540 308382 74592 308388
rect 70400 202156 70452 202162
rect 70400 202098 70452 202104
rect 69112 51740 69164 51746
rect 69112 51682 69164 51688
rect 69124 16574 69152 51682
rect 70412 16574 70440 202098
rect 73160 33788 73212 33794
rect 73160 33730 73212 33736
rect 73172 16574 73200 33730
rect 74552 16574 74580 308382
rect 81440 289128 81492 289134
rect 81440 289070 81492 289076
rect 77300 200796 77352 200802
rect 77300 200738 77352 200744
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72608 8968 72660 8974
rect 72608 8910 72660 8916
rect 72620 480 72648 8910
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 76196 9036 76248 9042
rect 76196 8978 76248 8984
rect 76208 480 76236 8978
rect 77312 3398 77340 200738
rect 81452 16574 81480 289070
rect 96620 279472 96672 279478
rect 96620 279414 96672 279420
rect 89720 278044 89772 278050
rect 89720 277986 89772 277992
rect 85580 276684 85632 276690
rect 85580 276626 85632 276632
rect 84200 214600 84252 214606
rect 84200 214542 84252 214548
rect 81452 16546 81664 16574
rect 80888 14544 80940 14550
rect 80888 14486 80940 14492
rect 77392 14476 77444 14482
rect 77392 14418 77444 14424
rect 77300 3392 77352 3398
rect 77300 3334 77352 3340
rect 77404 480 77432 14418
rect 79232 10328 79284 10334
rect 79232 10270 79284 10276
rect 78220 3392 78272 3398
rect 78220 3334 78272 3340
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78232 354 78260 3334
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 10270
rect 80900 480 80928 14486
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 10396 83332 10402
rect 83280 10338 83332 10344
rect 83292 480 83320 10338
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 214542
rect 85592 3398 85620 276626
rect 86960 213240 87012 213246
rect 86960 213182 87012 213188
rect 85672 35216 85724 35222
rect 85672 35158 85724 35164
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 85684 480 85712 35158
rect 86972 16574 87000 213182
rect 88340 199436 88392 199442
rect 88340 199378 88392 199384
rect 88352 16574 88380 199378
rect 89732 16574 89760 277986
rect 92480 198008 92532 198014
rect 92480 197950 92532 197956
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 14612 91612 14618
rect 91560 14554 91612 14560
rect 91572 480 91600 14554
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 197950
rect 95240 196648 95292 196654
rect 95240 196590 95292 196596
rect 95252 16574 95280 196590
rect 96632 16574 96660 279414
rect 100760 227044 100812 227050
rect 100760 226986 100812 226992
rect 98000 211812 98052 211818
rect 98000 211754 98052 211760
rect 98012 16574 98040 211754
rect 99380 62824 99432 62830
rect 99380 62766 99432 62772
rect 99392 16574 99420 62766
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93860 14680 93912 14686
rect 93860 14622 93912 14628
rect 93872 3398 93900 14622
rect 93952 13116 94004 13122
rect 93952 13058 94004 13064
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 13058
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 226986
rect 102152 3398 102180 336058
rect 103520 225616 103572 225622
rect 103520 225558 103572 225564
rect 102232 60036 102284 60042
rect 102232 59978 102284 59984
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 59978
rect 103532 16574 103560 225558
rect 104900 210452 104952 210458
rect 104900 210394 104952 210400
rect 104912 16574 104940 210394
rect 106280 195288 106332 195294
rect 106280 195230 106332 195236
rect 106292 16574 106320 195230
rect 110432 16574 110460 336126
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 110432 16546 110552 16574
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 109040 14748 109092 14754
rect 109040 14690 109092 14696
rect 108120 13184 108172 13190
rect 108120 13126 108172 13132
rect 108132 480 108160 13126
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 14690
rect 110524 480 110552 16546
rect 116400 15904 116452 15910
rect 116400 15846 116452 15852
rect 112352 14816 112404 14822
rect 112352 14758 112404 14764
rect 111616 13252 111668 13258
rect 111616 13194 111668 13200
rect 111628 480 111656 13194
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 14758
rect 114744 13320 114796 13326
rect 114744 13262 114796 13268
rect 114008 3324 114060 3330
rect 114008 3266 114060 3272
rect 114020 480 114048 3266
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 13262
rect 116412 480 116440 15846
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 336194
rect 224960 334688 225012 334694
rect 224960 334630 225012 334636
rect 175280 331968 175332 331974
rect 175280 331910 175332 331916
rect 168380 330608 168432 330614
rect 168380 330550 168432 330556
rect 164240 329180 164292 329186
rect 164240 329122 164292 329128
rect 125600 327752 125652 327758
rect 125600 327694 125652 327700
rect 118700 313948 118752 313954
rect 118700 313890 118752 313896
rect 118712 3398 118740 313890
rect 122840 311160 122892 311166
rect 122840 311102 122892 311108
rect 121460 280832 121512 280838
rect 121460 280774 121512 280780
rect 121472 16574 121500 280774
rect 122852 16574 122880 311102
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 118792 13388 118844 13394
rect 118792 13330 118844 13336
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 13330
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 121092 3324 121144 3330
rect 121092 3266 121144 3272
rect 121104 480 121132 3266
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 124692 480 124720 3198
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 327694
rect 160100 324964 160152 324970
rect 160100 324906 160152 324912
rect 128360 323672 128412 323678
rect 128360 323614 128412 323620
rect 126980 24132 127032 24138
rect 126980 24074 127032 24080
rect 126992 480 127020 24074
rect 128372 16574 128400 323614
rect 135260 309800 135312 309806
rect 135260 309742 135312 309748
rect 132500 308508 132552 308514
rect 132500 308450 132552 308456
rect 129740 273964 129792 273970
rect 129740 273906 129792 273912
rect 129752 16574 129780 273906
rect 131120 233912 131172 233918
rect 131120 233854 131172 233860
rect 131132 16574 131160 233854
rect 132512 16574 132540 308450
rect 133880 250504 133932 250510
rect 133880 250446 133932 250452
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128176 6180 128228 6186
rect 128176 6122 128228 6128
rect 128188 480 128216 6122
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 250446
rect 135272 4214 135300 309742
rect 146300 301504 146352 301510
rect 146300 301446 146352 301452
rect 143540 300144 143592 300150
rect 143540 300086 143592 300092
rect 136640 290488 136692 290494
rect 136640 290430 136692 290436
rect 135352 54528 135404 54534
rect 135352 54470 135404 54476
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 135364 3482 135392 54470
rect 136652 16574 136680 290430
rect 139400 287700 139452 287706
rect 139400 287642 139452 287648
rect 138020 36576 138072 36582
rect 138020 36518 138072 36524
rect 138032 16574 138060 36518
rect 139412 16574 139440 287642
rect 140780 247716 140832 247722
rect 140780 247658 140832 247664
rect 140792 16574 140820 247658
rect 142160 228404 142212 228410
rect 142160 228346 142212 228352
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 4150
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 228346
rect 143552 480 143580 300086
rect 143632 246356 143684 246362
rect 143632 246298 143684 246304
rect 143644 16574 143672 246298
rect 144920 21412 144972 21418
rect 144920 21354 144972 21360
rect 144932 16574 144960 21354
rect 146312 16574 146340 301446
rect 154580 291848 154632 291854
rect 154580 291790 154632 291796
rect 150440 272536 150492 272542
rect 150440 272478 150492 272484
rect 147680 244928 147732 244934
rect 147680 244870 147732 244876
rect 147692 16574 147720 244870
rect 149060 53100 149112 53106
rect 149060 53042 149112 53048
rect 149072 16574 149100 53042
rect 150452 16574 150480 272478
rect 153200 271176 153252 271182
rect 153200 271118 153252 271124
rect 151820 243568 151872 243574
rect 151820 243510 151872 243516
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 243510
rect 151912 55888 151964 55894
rect 151912 55830 151964 55836
rect 151924 16574 151952 55830
rect 153212 16574 153240 271118
rect 154592 16574 154620 291790
rect 157340 289196 157392 289202
rect 157340 289138 157392 289144
rect 155960 57248 156012 57254
rect 155960 57190 156012 57196
rect 155972 16574 156000 57190
rect 157352 16574 157380 289138
rect 158720 242208 158772 242214
rect 158720 242150 158772 242156
rect 158732 16574 158760 242150
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11830 160140 324906
rect 161480 269816 161532 269822
rect 161480 269758 161532 269764
rect 160192 58676 160244 58682
rect 160192 58618 160244 58624
rect 160100 11824 160152 11830
rect 160100 11766 160152 11772
rect 160204 6914 160232 58618
rect 161492 16574 161520 269758
rect 162860 25628 162912 25634
rect 162860 25570 162912 25576
rect 162872 16574 162900 25570
rect 164252 16574 164280 329122
rect 165620 268388 165672 268394
rect 165620 268330 165672 268336
rect 165632 16574 165660 268330
rect 167000 239420 167052 239426
rect 167000 239362 167052 239368
rect 167012 16574 167040 239362
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 11824 161348 11830
rect 161296 11766 161348 11772
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11766
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 330550
rect 171140 312656 171192 312662
rect 171140 312598 171192 312604
rect 168472 265668 168524 265674
rect 168472 265610 168524 265616
rect 168484 16574 168512 265610
rect 169760 37936 169812 37942
rect 169760 37878 169812 37884
rect 169772 16574 169800 37878
rect 171152 16574 171180 312598
rect 172520 264240 172572 264246
rect 172520 264182 172572 264188
rect 172532 16574 172560 264182
rect 175292 16574 175320 331910
rect 201500 327820 201552 327826
rect 201500 327762 201552 327768
rect 193220 326460 193272 326466
rect 193220 326402 193272 326408
rect 176660 325032 176712 325038
rect 176660 324974 176712 324980
rect 168484 16546 169616 16574
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 175292 16546 175504 16574
rect 169588 480 169616 16546
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173900 10464 173952 10470
rect 173900 10406 173952 10412
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 10406
rect 175476 480 175504 16546
rect 176672 4214 176700 324974
rect 189080 322312 189132 322318
rect 189080 322254 189132 322260
rect 179420 303000 179472 303006
rect 179420 302942 179472 302948
rect 178040 286408 178092 286414
rect 178040 286350 178092 286356
rect 178052 16574 178080 286350
rect 179432 16574 179460 302942
rect 182180 285048 182232 285054
rect 182180 284990 182232 284996
rect 180800 238060 180852 238066
rect 180800 238002 180852 238008
rect 180812 16574 180840 238002
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 176752 7608 176804 7614
rect 176752 7550 176804 7556
rect 176660 4208 176712 4214
rect 176660 4150 176712 4156
rect 176764 3482 176792 7550
rect 177856 4208 177908 4214
rect 177856 4150 177908 4156
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 4150
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 284990
rect 184940 283688 184992 283694
rect 184940 283630 184992 283636
rect 183560 262880 183612 262886
rect 183560 262822 183612 262828
rect 183572 16574 183600 262822
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 283630
rect 186320 261520 186372 261526
rect 186320 261462 186372 261468
rect 185032 39364 185084 39370
rect 185032 39306 185084 39312
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 185044 6914 185072 39306
rect 186332 16574 186360 261462
rect 187700 236700 187752 236706
rect 187700 236642 187752 236648
rect 187712 16574 187740 236642
rect 189092 16574 189120 322254
rect 190460 260160 190512 260166
rect 190460 260102 190512 260108
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 260102
rect 191840 235272 191892 235278
rect 191840 235214 191892 235220
rect 191852 16574 191880 235214
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 326402
rect 195980 282260 196032 282266
rect 195980 282202 196032 282208
rect 193312 258800 193364 258806
rect 193312 258742 193364 258748
rect 193324 16574 193352 258742
rect 194600 40724 194652 40730
rect 194600 40666 194652 40672
rect 194612 16574 194640 40666
rect 195992 16574 196020 282202
rect 200120 280900 200172 280906
rect 200120 280842 200172 280848
rect 198740 42084 198792 42090
rect 198740 42026 198792 42032
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197912 7676 197964 7682
rect 197912 7618 197964 7624
rect 197924 480 197952 7618
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 42026
rect 200132 16574 200160 280842
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 327762
rect 215300 320884 215352 320890
rect 215300 320826 215352 320832
rect 205640 319456 205692 319462
rect 205640 319398 205692 319404
rect 202880 279540 202932 279546
rect 202880 279482 202932 279488
rect 201592 232552 201644 232558
rect 201592 232494 201644 232500
rect 201604 16574 201632 232494
rect 202892 16574 202920 279482
rect 204260 257440 204312 257446
rect 204260 257382 204312 257388
rect 204272 16574 204300 257382
rect 205652 16574 205680 319398
rect 207020 307148 207072 307154
rect 207020 307090 207072 307096
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 307090
rect 209780 304360 209832 304366
rect 209780 304302 209832 304308
rect 208400 256080 208452 256086
rect 208400 256022 208452 256028
rect 208412 16574 208440 256022
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 9674 209820 304302
rect 213920 278112 213972 278118
rect 213920 278054 213972 278060
rect 211160 254652 211212 254658
rect 211160 254594 211212 254600
rect 209872 231124 209924 231130
rect 209872 231066 209924 231072
rect 209700 9654 209820 9674
rect 209688 9648 209820 9654
rect 209740 9646 209820 9648
rect 209688 9590 209740 9596
rect 209884 6914 209912 231066
rect 211172 16574 211200 254594
rect 212540 229764 212592 229770
rect 212540 229706 212592 229712
rect 212552 16574 212580 229706
rect 213932 16574 213960 278054
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 9648 211028 9654
rect 210976 9590 211028 9596
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 210988 480 211016 9590
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 320826
rect 219440 318096 219492 318102
rect 219440 318038 219492 318044
rect 216680 43444 216732 43450
rect 216680 43386 216732 43392
rect 216692 16574 216720 43386
rect 218060 26920 218112 26926
rect 218060 26862 218112 26868
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 3194 218100 26862
rect 219452 16574 219480 318038
rect 223580 316736 223632 316742
rect 223580 316678 223632 316684
rect 220820 276752 220872 276758
rect 220820 276694 220872 276700
rect 220832 16574 220860 276694
rect 222200 267028 222252 267034
rect 222200 266970 222252 266976
rect 222212 16574 222240 266970
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 218152 4820 218204 4826
rect 218152 4762 218204 4768
rect 218060 3188 218112 3194
rect 218060 3130 218112 3136
rect 218164 2394 218192 4762
rect 219256 3188 219308 3194
rect 219256 3130 219308 3136
rect 218072 2366 218192 2394
rect 218072 480 218100 2366
rect 219268 480 219296 3130
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 316678
rect 224972 16574 225000 334630
rect 226340 315308 226392 315314
rect 226340 315250 226392 315256
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 11830 226380 315250
rect 227720 275392 227772 275398
rect 227720 275334 227772 275340
rect 226432 253292 226484 253298
rect 226432 253234 226484 253240
rect 226340 11824 226392 11830
rect 226340 11766 226392 11772
rect 226444 6914 226472 253234
rect 227732 16574 227760 275334
rect 227732 16546 228312 16574
rect 227536 11824 227588 11830
rect 227536 11766 227588 11772
rect 226352 6886 226472 6914
rect 226352 480 226380 6886
rect 227548 480 227576 11766
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228376 4826 228404 336262
rect 229100 251932 229152 251938
rect 229100 251874 229152 251880
rect 229112 16574 229140 251874
rect 229756 164218 229784 460974
rect 233884 458788 233936 458794
rect 233884 458730 233936 458736
rect 232504 458652 232556 458658
rect 232504 458594 232556 458600
rect 231216 458584 231268 458590
rect 231216 458526 231268 458532
rect 231124 336388 231176 336394
rect 231124 336330 231176 336336
rect 229744 164212 229796 164218
rect 229744 164154 229796 164160
rect 230480 44872 230532 44878
rect 230480 44814 230532 44820
rect 230492 16574 230520 44814
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 228364 4820 228416 4826
rect 228364 4762 228416 4768
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 231136 6186 231164 336330
rect 231228 267714 231256 458526
rect 231860 333192 231912 333198
rect 231860 333134 231912 333140
rect 231216 267708 231268 267714
rect 231216 267650 231268 267656
rect 231124 6180 231176 6186
rect 231124 6122 231176 6128
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 333134
rect 232516 320142 232544 458594
rect 233896 372570 233924 458730
rect 233988 449886 234016 461314
rect 266372 460154 266400 697546
rect 298100 643136 298152 643142
rect 298100 643078 298152 643084
rect 296720 616888 296772 616894
rect 296720 616830 296772 616836
rect 293960 590708 294012 590714
rect 293960 590650 294012 590656
rect 292580 563100 292632 563106
rect 292580 563042 292632 563048
rect 288440 536852 288492 536858
rect 288440 536794 288492 536800
rect 287060 510672 287112 510678
rect 287060 510614 287112 510620
rect 284300 484424 284352 484430
rect 284300 484366 284352 484372
rect 277124 462460 277176 462466
rect 277124 462402 277176 462408
rect 273996 461168 274048 461174
rect 273996 461110 274048 461116
rect 266360 460148 266412 460154
rect 266360 460090 266412 460096
rect 255044 458516 255096 458522
rect 255044 458458 255096 458464
rect 245568 458448 245620 458454
rect 245568 458390 245620 458396
rect 240784 458380 240836 458386
rect 240784 458322 240836 458328
rect 235908 458312 235960 458318
rect 235908 458254 235960 458260
rect 235920 457994 235948 458254
rect 240796 457994 240824 458322
rect 245580 457994 245608 458390
rect 255056 457994 255084 458458
rect 274008 457994 274036 461110
rect 275560 458720 275612 458726
rect 275560 458662 275612 458668
rect 275572 457994 275600 458662
rect 277136 457994 277164 462402
rect 280068 461304 280120 461310
rect 280068 461246 280120 461252
rect 278688 461236 278740 461242
rect 278688 461178 278740 461184
rect 278700 457994 278728 461178
rect 280080 457994 280108 461246
rect 235796 457966 235948 457994
rect 240488 457966 240824 457994
rect 245272 457966 245608 457994
rect 254748 457966 255084 457994
rect 273700 457966 274036 457994
rect 275264 457966 275600 457994
rect 276828 457966 277164 457994
rect 278392 457966 278728 457994
rect 279956 457966 280108 457994
rect 284312 457994 284340 484366
rect 287072 480254 287100 510614
rect 288452 480254 288480 536794
rect 289820 524476 289872 524482
rect 289820 524418 289872 524424
rect 289832 480254 289860 524418
rect 287072 480226 287468 480254
rect 288452 480226 289032 480254
rect 289832 480226 290596 480254
rect 285864 470620 285916 470626
rect 285864 470562 285916 470568
rect 285876 457994 285904 470562
rect 287440 457994 287468 480226
rect 289004 457994 289032 480226
rect 290568 457994 290596 480226
rect 292592 457994 292620 563042
rect 293972 457994 294000 590650
rect 295340 576904 295392 576910
rect 295340 576846 295392 576852
rect 295352 457994 295380 576846
rect 296732 480254 296760 616830
rect 298112 480254 298140 643078
rect 296732 480226 296944 480254
rect 298112 480226 298508 480254
rect 296916 457994 296944 480226
rect 298480 457994 298508 480226
rect 299492 467158 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 328460 700868 328512 700874
rect 328460 700810 328512 700816
rect 318800 700800 318852 700806
rect 318800 700742 318852 700748
rect 314660 700664 314712 700670
rect 314660 700606 314712 700612
rect 303620 696992 303672 696998
rect 303620 696934 303672 696940
rect 300860 670812 300912 670818
rect 300860 670754 300912 670760
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299584 480254 299612 630634
rect 300872 480254 300900 670754
rect 299584 480226 300072 480254
rect 300872 480226 301728 480254
rect 299480 467152 299532 467158
rect 299480 467094 299532 467100
rect 300044 457994 300072 480226
rect 301700 457994 301728 480226
rect 303632 457994 303660 696934
rect 305000 683188 305052 683194
rect 305000 683130 305052 683136
rect 305012 457994 305040 683130
rect 311164 464364 311216 464370
rect 311164 464306 311216 464312
rect 307116 461644 307168 461650
rect 307116 461586 307168 461592
rect 307128 457994 307156 461586
rect 308680 460624 308732 460630
rect 308680 460566 308732 460572
rect 308692 457994 308720 460566
rect 310244 460556 310296 460562
rect 310244 460498 310296 460504
rect 310256 457994 310284 460498
rect 284312 457966 284740 457994
rect 285876 457966 286304 457994
rect 287440 457966 287868 457994
rect 289004 457966 289432 457994
rect 290568 457966 290996 457994
rect 292592 457966 292652 457994
rect 293972 457966 294216 457994
rect 295352 457966 295780 457994
rect 296916 457966 297344 457994
rect 298480 457966 298908 457994
rect 300044 457966 300472 457994
rect 301700 457966 302128 457994
rect 303632 457966 303692 457994
rect 305012 457966 305256 457994
rect 306820 457966 307156 457994
rect 308384 457966 308720 457994
rect 309948 457966 310284 457994
rect 311176 457994 311204 464306
rect 313096 460760 313148 460766
rect 313096 460702 313148 460708
rect 311176 457966 311604 457994
rect 313108 457858 313136 460702
rect 314672 457994 314700 700606
rect 318812 480254 318840 700742
rect 320180 502988 320232 502994
rect 320180 502930 320232 502936
rect 320192 480254 320220 502930
rect 318812 480226 319024 480254
rect 320192 480226 320680 480254
rect 316040 465724 316092 465730
rect 316040 465666 316092 465672
rect 316052 457994 316080 465666
rect 318156 460896 318208 460902
rect 318156 460838 318208 460844
rect 318168 457994 318196 460838
rect 314672 457966 314732 457994
rect 316052 457966 316296 457994
rect 317860 457966 318196 457994
rect 318996 457994 319024 480226
rect 320652 457994 320680 480226
rect 325700 467152 325752 467158
rect 325700 467094 325752 467100
rect 324136 460080 324188 460086
rect 324136 460022 324188 460028
rect 322848 460012 322900 460018
rect 322848 459954 322900 459960
rect 322860 457994 322888 459954
rect 318996 457966 319424 457994
rect 320652 457966 321080 457994
rect 322644 457966 322888 457994
rect 324148 457858 324176 460022
rect 325712 457994 325740 467094
rect 327080 460148 327132 460154
rect 327080 460090 327132 460096
rect 327092 457994 327120 460090
rect 328472 457994 328500 700810
rect 329840 698964 329892 698970
rect 329840 698906 329892 698912
rect 329852 480254 329880 698906
rect 329852 480226 330156 480254
rect 330128 457994 330156 480226
rect 331232 460018 331260 702986
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332600 700732 332652 700738
rect 332600 700674 332652 700680
rect 332612 480254 332640 700674
rect 338120 700596 338172 700602
rect 338120 700538 338172 700544
rect 332612 480226 333284 480254
rect 331772 460828 331824 460834
rect 331772 460770 331824 460776
rect 331220 460012 331272 460018
rect 331220 459954 331272 459960
rect 331784 457994 331812 460770
rect 333256 457994 333284 480226
rect 334808 468512 334860 468518
rect 334808 468454 334860 468460
rect 334820 457994 334848 468454
rect 336740 460692 336792 460698
rect 336740 460634 336792 460640
rect 336752 457994 336780 460634
rect 338132 457994 338160 700538
rect 342260 700528 342312 700534
rect 342260 700470 342312 700476
rect 340880 700460 340932 700466
rect 340880 700402 340932 700408
rect 340892 480254 340920 700402
rect 342272 480254 342300 700470
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 345032 480254 345060 700266
rect 340892 480226 341196 480254
rect 342272 480226 342760 480254
rect 345032 480226 345888 480254
rect 339684 460488 339736 460494
rect 339684 460430 339736 460436
rect 339696 457994 339724 460430
rect 341168 457994 341196 480226
rect 342732 457994 342760 480226
rect 344374 460320 344430 460329
rect 344374 460255 344430 460264
rect 344388 457994 344416 460255
rect 345860 457994 345888 480226
rect 347792 460086 347820 702406
rect 347872 700392 347924 700398
rect 347872 700334 347924 700340
rect 347780 460080 347832 460086
rect 347780 460022 347832 460028
rect 347884 458266 347912 700334
rect 351920 670744 351972 670750
rect 351920 670686 351972 670692
rect 350540 656940 350592 656946
rect 350540 656882 350592 656888
rect 350552 480254 350580 656882
rect 351932 480254 351960 670686
rect 356060 618316 356112 618322
rect 356060 618258 356112 618264
rect 354680 605872 354732 605878
rect 354680 605814 354732 605820
rect 354692 480254 354720 605814
rect 356072 480254 356100 618258
rect 361580 565888 361632 565894
rect 361580 565830 361632 565836
rect 360200 553444 360252 553450
rect 360200 553386 360252 553392
rect 350552 480226 350672 480254
rect 351932 480226 352236 480254
rect 354692 480226 355364 480254
rect 356072 480226 356928 480254
rect 349158 460184 349214 460193
rect 349158 460119 349214 460128
rect 349068 459604 349120 459610
rect 349068 459546 349120 459552
rect 349080 458862 349108 459546
rect 349068 458856 349120 458862
rect 349068 458798 349120 458804
rect 347838 458238 347912 458266
rect 325712 457966 325772 457994
rect 327092 457966 327336 457994
rect 328472 457966 328900 457994
rect 330128 457966 330556 457994
rect 331784 457966 332120 457994
rect 333256 457966 333684 457994
rect 334820 457966 335248 457994
rect 336752 457966 336812 457994
rect 338132 457966 338376 457994
rect 339696 457966 340032 457994
rect 341168 457966 341596 457994
rect 342732 457966 343160 457994
rect 344388 457966 344724 457994
rect 345860 457966 346288 457994
rect 347838 457980 347866 458238
rect 349172 457994 349200 460119
rect 349804 459672 349856 459678
rect 349804 459614 349856 459620
rect 349172 457966 349508 457994
rect 313108 457830 313168 457858
rect 324148 457830 324208 457858
rect 281632 457632 281684 457638
rect 281520 457580 281632 457586
rect 281520 457574 281684 457580
rect 281520 457558 281672 457574
rect 349816 457502 349844 459614
rect 350644 457994 350672 480226
rect 352208 457994 352236 480226
rect 353852 460420 353904 460426
rect 353852 460362 353904 460368
rect 353864 457994 353892 460362
rect 355336 457994 355364 480226
rect 356900 457994 356928 480226
rect 358820 460352 358872 460358
rect 358820 460294 358872 460300
rect 358832 457994 358860 460294
rect 360212 457994 360240 553386
rect 361592 480254 361620 565830
rect 364352 502994 364380 702406
rect 365720 514820 365772 514826
rect 365720 514762 365772 514768
rect 364340 502988 364392 502994
rect 364340 502930 364392 502936
rect 364340 501016 364392 501022
rect 364340 500958 364392 500964
rect 364352 480254 364380 500958
rect 365732 480254 365760 514762
rect 361592 480226 361712 480254
rect 364352 480226 364840 480254
rect 365732 480226 366404 480254
rect 361684 457994 361712 480226
rect 363328 460284 363380 460290
rect 363328 460226 363380 460232
rect 363340 457994 363368 460226
rect 364812 457994 364840 480226
rect 366376 457994 366404 480226
rect 375932 462528 375984 462534
rect 375932 462470 375984 462476
rect 371240 462392 371292 462398
rect 371240 462334 371292 462340
rect 369860 461372 369912 461378
rect 369860 461314 369912 461320
rect 368112 460216 368164 460222
rect 368112 460158 368164 460164
rect 368124 457994 368152 460158
rect 369872 457994 369900 461314
rect 371252 457994 371280 462334
rect 374368 459672 374420 459678
rect 374368 459614 374420 459620
rect 373126 458244 373178 458250
rect 373126 458186 373178 458192
rect 350644 457966 351072 457994
rect 352208 457966 352636 457994
rect 353864 457966 354200 457994
rect 355336 457966 355764 457994
rect 356900 457966 357328 457994
rect 358832 457966 358984 457994
rect 360212 457966 360548 457994
rect 361684 457966 362112 457994
rect 363340 457966 363676 457994
rect 364812 457966 365240 457994
rect 366376 457966 366804 457994
rect 368124 457966 368460 457994
rect 369872 457966 370024 457994
rect 371252 457966 371588 457994
rect 373138 457980 373166 458186
rect 374380 457994 374408 459614
rect 375944 457994 375972 462470
rect 379152 461100 379204 461106
rect 379152 461042 379204 461048
rect 377588 458788 377640 458794
rect 377588 458730 377640 458736
rect 377600 457994 377628 458730
rect 379164 457994 379192 461042
rect 396540 461032 396592 461038
rect 396540 460974 396592 460980
rect 391940 460964 391992 460970
rect 391940 460906 391992 460912
rect 380900 459604 380952 459610
rect 380900 459546 380952 459552
rect 380912 457994 380940 459546
rect 382280 458652 382332 458658
rect 382280 458594 382332 458600
rect 382292 457994 382320 458594
rect 387064 458584 387116 458590
rect 387064 458526 387116 458532
rect 387076 457994 387104 458526
rect 391952 457994 391980 460906
rect 396552 457994 396580 460974
rect 397472 460902 397500 703520
rect 413664 700806 413692 703520
rect 413652 700800 413704 700806
rect 413652 700742 413704 700748
rect 429212 465730 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 465724 429252 465730
rect 429200 465666 429252 465672
rect 425704 462460 425756 462466
rect 425704 462402 425756 462408
rect 417516 461304 417568 461310
rect 417516 461246 417568 461252
rect 397460 460896 397512 460902
rect 397460 460838 397512 460844
rect 407578 459776 407634 459785
rect 407578 459711 407634 459720
rect 407592 457994 407620 459711
rect 417424 458380 417476 458386
rect 417424 458322 417476 458328
rect 374380 457966 374716 457994
rect 375944 457966 376280 457994
rect 377600 457966 377936 457994
rect 379164 457966 379500 457994
rect 380912 457966 381064 457994
rect 382292 457966 382628 457994
rect 387076 457966 387412 457994
rect 391952 457966 392104 457994
rect 396552 457966 396888 457994
rect 407592 457966 407928 457994
rect 283380 457496 283432 457502
rect 237654 457464 237710 457473
rect 237360 457422 237654 457450
rect 239218 457464 239274 457473
rect 238924 457422 239218 457450
rect 237654 457399 237710 457408
rect 242346 457464 242402 457473
rect 242052 457422 242346 457450
rect 239218 457399 239274 457408
rect 243910 457464 243966 457473
rect 243616 457422 243910 457450
rect 242346 457399 242402 457408
rect 243910 457399 243966 457408
rect 246670 457464 246726 457473
rect 248234 457464 248290 457473
rect 246726 457422 246836 457450
rect 246670 457399 246726 457408
rect 250258 457464 250314 457473
rect 248290 457422 248400 457450
rect 249964 457422 250258 457450
rect 248234 457399 248290 457408
rect 251822 457464 251878 457473
rect 251528 457422 251822 457450
rect 250258 457399 250314 457408
rect 253386 457464 253442 457473
rect 253092 457422 253386 457450
rect 251822 457399 251878 457408
rect 256514 457464 256570 457473
rect 256312 457422 256514 457450
rect 253386 457399 253442 457408
rect 256514 457399 256570 457408
rect 257710 457464 257766 457473
rect 259274 457464 259330 457473
rect 257766 457422 257876 457450
rect 257710 457399 257766 457408
rect 261298 457464 261354 457473
rect 259330 457422 259440 457450
rect 261004 457422 261298 457450
rect 259274 457399 259330 457408
rect 262862 457464 262918 457473
rect 262568 457422 262862 457450
rect 261298 457399 261354 457408
rect 264518 457464 264574 457473
rect 264224 457422 264518 457450
rect 262862 457399 262918 457408
rect 266082 457464 266138 457473
rect 265788 457422 266082 457450
rect 264518 457399 264574 457408
rect 267554 457464 267610 457473
rect 267352 457422 267554 457450
rect 266082 457399 266138 457408
rect 267554 457399 267610 457408
rect 268750 457464 268806 457473
rect 270590 457464 270646 457473
rect 268806 457422 268916 457450
rect 270480 457422 270590 457450
rect 268750 457399 268806 457408
rect 272338 457464 272394 457473
rect 272044 457422 272338 457450
rect 270590 457399 270646 457408
rect 283176 457444 283380 457450
rect 283176 457438 283432 457444
rect 349804 457496 349856 457502
rect 349804 457438 349856 457444
rect 383842 457464 383898 457473
rect 283176 457422 283420 457438
rect 272338 457399 272394 457408
rect 385406 457464 385462 457473
rect 383898 457422 384192 457450
rect 383842 457399 383898 457408
rect 388626 457464 388682 457473
rect 385462 457422 385756 457450
rect 385406 457399 385462 457408
rect 390190 457464 390246 457473
rect 388682 457422 388976 457450
rect 388626 457399 388682 457408
rect 393502 457464 393558 457473
rect 390246 457422 390540 457450
rect 390190 457399 390246 457408
rect 394882 457464 394938 457473
rect 393558 457422 393668 457450
rect 393502 457399 393558 457408
rect 398102 457464 398158 457473
rect 394938 457422 395232 457450
rect 394882 457399 394938 457408
rect 399666 457464 399722 457473
rect 398158 457422 398452 457450
rect 398102 457399 398158 457408
rect 401230 457464 401286 457473
rect 399722 457422 400016 457450
rect 399666 457399 399722 457408
rect 402978 457464 403034 457473
rect 401286 457422 401580 457450
rect 401230 457399 401286 457408
rect 404358 457464 404414 457473
rect 403034 457422 403144 457450
rect 402978 457399 403034 457408
rect 406014 457464 406070 457473
rect 404414 457422 404708 457450
rect 404358 457399 404414 457408
rect 409142 457464 409198 457473
rect 406070 457422 406364 457450
rect 406014 457399 406070 457408
rect 410706 457464 410762 457473
rect 409198 457422 409492 457450
rect 409142 457399 409198 457408
rect 412270 457464 412326 457473
rect 410762 457422 411056 457450
rect 410706 457399 410762 457408
rect 412326 457422 412620 457450
rect 414184 457422 414980 457450
rect 412270 457399 412326 457408
rect 233976 449880 234028 449886
rect 233976 449822 234028 449828
rect 233884 372564 233936 372570
rect 233884 372506 233936 372512
rect 270696 338150 270940 338178
rect 234816 338014 235152 338042
rect 235276 338014 235428 338042
rect 235552 338014 235796 338042
rect 236104 338014 236164 338042
rect 236288 338014 236532 338042
rect 236656 338014 236900 338042
rect 237024 338014 237268 338042
rect 237576 338014 237636 338042
rect 237760 338014 238004 338042
rect 238128 338014 238372 338042
rect 238496 338014 238740 338042
rect 238864 338014 239108 338042
rect 239232 338014 239476 338042
rect 239600 338014 239844 338042
rect 240152 338014 240212 338042
rect 240336 338014 240580 338042
rect 240704 338014 240948 338042
rect 241072 338014 241316 338042
rect 241684 338014 241836 338042
rect 233976 335368 234028 335374
rect 233976 335310 234028 335316
rect 233882 334656 233938 334665
rect 233882 334591 233938 334600
rect 232504 320136 232556 320142
rect 232504 320078 232556 320084
rect 232594 319424 232650 319433
rect 232594 319359 232650 319368
rect 232608 241466 232636 319359
rect 233240 249144 233292 249150
rect 233240 249086 233292 249092
rect 232596 241460 232648 241466
rect 232596 241402 232648 241408
rect 233252 16574 233280 249086
rect 233896 71738 233924 334591
rect 233988 249082 234016 335310
rect 234816 334626 234844 338014
rect 235276 335354 235304 338014
rect 234908 335326 235304 335354
rect 234804 334620 234856 334626
rect 234804 334562 234856 334568
rect 234908 321554 234936 335326
rect 234724 321526 234936 321554
rect 234724 275330 234752 321526
rect 235552 316034 235580 338014
rect 234816 316006 235580 316034
rect 234712 275324 234764 275330
rect 234712 275266 234764 275272
rect 233976 249076 234028 249082
rect 233976 249018 234028 249024
rect 234816 111110 234844 316006
rect 236104 286346 236132 338014
rect 236092 286340 236144 286346
rect 236092 286282 236144 286288
rect 234804 111104 234856 111110
rect 234804 111046 234856 111052
rect 233884 71732 233936 71738
rect 233884 71674 233936 71680
rect 234620 46232 234672 46238
rect 234620 46174 234672 46180
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 480 234660 46174
rect 235816 6316 235868 6322
rect 235816 6258 235868 6264
rect 235828 480 235856 6258
rect 236288 3369 236316 338014
rect 236656 336054 236684 338014
rect 236644 336048 236696 336054
rect 236644 335990 236696 335996
rect 237024 326398 237052 338014
rect 237576 326534 237604 338014
rect 237760 335354 237788 338014
rect 237668 335326 237788 335354
rect 237564 326528 237616 326534
rect 237564 326470 237616 326476
rect 237012 326392 237064 326398
rect 237012 326334 237064 326340
rect 237380 326392 237432 326398
rect 237380 326334 237432 326340
rect 237012 6248 237064 6254
rect 237012 6190 237064 6196
rect 236274 3360 236330 3369
rect 236274 3295 236330 3304
rect 237024 480 237052 6190
rect 237392 3505 237420 326334
rect 237668 321586 237696 335326
rect 237748 326528 237800 326534
rect 237748 326470 237800 326476
rect 237484 321558 237696 321586
rect 237484 97306 237512 321558
rect 237760 318794 237788 326470
rect 238128 326398 238156 338014
rect 238116 326392 238168 326398
rect 238116 326334 238168 326340
rect 237576 318766 237788 318794
rect 237576 222902 237604 318766
rect 238496 316034 238524 338014
rect 238760 326392 238812 326398
rect 238760 326334 238812 326340
rect 237668 316006 238524 316034
rect 237668 302938 237696 316006
rect 237656 302932 237708 302938
rect 237656 302874 237708 302880
rect 237564 222896 237616 222902
rect 237564 222838 237616 222844
rect 237472 97300 237524 97306
rect 237472 97242 237524 97248
rect 237472 47592 237524 47598
rect 237472 47534 237524 47540
rect 237484 16574 237512 47534
rect 237484 16546 237696 16574
rect 237378 3496 237434 3505
rect 237378 3431 237434 3440
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 354 237696 16546
rect 238772 3466 238800 326334
rect 238864 11762 238892 338014
rect 239232 316034 239260 338014
rect 239600 326398 239628 338014
rect 240152 335374 240180 338014
rect 240140 335368 240192 335374
rect 240140 335310 240192 335316
rect 239588 326392 239640 326398
rect 239588 326334 239640 326340
rect 240232 326392 240284 326398
rect 240232 326334 240284 326340
rect 238956 316006 239260 316034
rect 238956 258738 238984 316006
rect 238944 258732 238996 258738
rect 238944 258674 238996 258680
rect 238852 11756 238904 11762
rect 238852 11698 238904 11704
rect 239312 11756 239364 11762
rect 239312 11698 239364 11704
rect 238760 3460 238812 3466
rect 238760 3402 238812 3408
rect 239324 480 239352 11698
rect 240244 3602 240272 326334
rect 240336 256018 240364 338014
rect 240704 326398 240732 338014
rect 240692 326392 240744 326398
rect 240692 326334 240744 326340
rect 241072 316034 241100 338014
rect 241808 326534 241836 338014
rect 241900 338014 242052 338042
rect 242176 338014 242420 338042
rect 242544 338014 242788 338042
rect 241796 326528 241848 326534
rect 241796 326470 241848 326476
rect 241612 326392 241664 326398
rect 241612 326334 241664 326340
rect 241520 326324 241572 326330
rect 241520 326266 241572 326272
rect 240428 316006 241100 316034
rect 240324 256012 240376 256018
rect 240324 255954 240376 255960
rect 240324 28280 240376 28286
rect 240324 28222 240376 28228
rect 240232 3596 240284 3602
rect 240232 3538 240284 3544
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240336 354 240364 28222
rect 240428 3534 240456 316006
rect 241532 3738 241560 326266
rect 241520 3732 241572 3738
rect 241520 3674 241572 3680
rect 241624 3670 241652 326334
rect 241900 323626 241928 338014
rect 241980 326528 242032 326534
rect 241980 326470 242032 326476
rect 241716 323598 241928 323626
rect 241716 257378 241744 323598
rect 241992 318794 242020 326470
rect 242176 326398 242204 338014
rect 242164 326392 242216 326398
rect 242164 326334 242216 326340
rect 242544 326330 242572 338014
rect 243142 337770 243170 338028
rect 243280 338014 243524 338042
rect 243648 338014 243892 338042
rect 244016 338014 244260 338042
rect 244384 338014 244628 338042
rect 244752 338014 244996 338042
rect 245120 338014 245364 338042
rect 245732 338014 245884 338042
rect 243142 337742 243216 337770
rect 242992 336728 243044 336734
rect 242992 336670 243044 336676
rect 242532 326324 242584 326330
rect 242532 326266 242584 326272
rect 242900 326052 242952 326058
rect 242900 325994 242952 326000
rect 241808 318766 242020 318794
rect 241808 282198 241836 318766
rect 241796 282192 241848 282198
rect 241796 282134 241848 282140
rect 241704 257372 241756 257378
rect 241704 257314 241756 257320
rect 241704 17264 241756 17270
rect 241704 17206 241756 17212
rect 241612 3664 241664 3670
rect 241612 3606 241664 3612
rect 240416 3528 240468 3534
rect 240416 3470 240468 3476
rect 241716 480 241744 17206
rect 242912 3806 242940 325994
rect 243004 68338 243032 336670
rect 243188 323610 243216 337742
rect 243280 336734 243308 338014
rect 243268 336728 243320 336734
rect 243268 336670 243320 336676
rect 243648 326058 243676 338014
rect 243636 326052 243688 326058
rect 243636 325994 243688 326000
rect 243176 323604 243228 323610
rect 243176 323546 243228 323552
rect 244016 321554 244044 338014
rect 244280 330472 244332 330478
rect 244280 330414 244332 330420
rect 243096 321526 244044 321554
rect 243096 251870 243124 321526
rect 243084 251864 243136 251870
rect 243084 251806 243136 251812
rect 242992 68332 243044 68338
rect 242992 68274 243044 68280
rect 242992 29640 243044 29646
rect 242992 29582 243044 29588
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 242900 3596 242952 3602
rect 242900 3538 242952 3544
rect 242912 480 242940 3538
rect 243004 3482 243032 29582
rect 243084 17332 243136 17338
rect 243084 17274 243136 17280
rect 243096 3602 243124 17274
rect 244292 3874 244320 330414
rect 244384 209098 244412 338014
rect 244752 330478 244780 338014
rect 245120 336682 245148 338014
rect 244844 336654 245148 336682
rect 244740 330472 244792 330478
rect 244740 330414 244792 330420
rect 244844 316034 244872 336654
rect 244924 336592 244976 336598
rect 244924 336534 244976 336540
rect 244476 316006 244872 316034
rect 244476 253230 244504 316006
rect 244936 283626 244964 336534
rect 245752 328568 245804 328574
rect 245752 328510 245804 328516
rect 244924 283620 244976 283626
rect 244924 283562 244976 283568
rect 244464 253224 244516 253230
rect 244464 253166 244516 253172
rect 244372 209092 244424 209098
rect 244372 209034 244424 209040
rect 244372 49020 244424 49026
rect 244372 48962 244424 48968
rect 244384 16574 244412 48962
rect 245764 18630 245792 328510
rect 245856 254590 245884 338014
rect 245948 338014 246100 338042
rect 246224 338014 246468 338042
rect 246592 338014 246836 338042
rect 245844 254584 245896 254590
rect 245844 254526 245896 254532
rect 245752 18624 245804 18630
rect 245752 18566 245804 18572
rect 244384 16546 245240 16574
rect 244280 3868 244332 3874
rect 244280 3810 244332 3816
rect 243084 3596 243136 3602
rect 243084 3538 243136 3544
rect 243004 3454 244136 3482
rect 244108 480 244136 3454
rect 245212 480 245240 16546
rect 245948 3942 245976 338014
rect 246224 336598 246252 338014
rect 246304 336728 246356 336734
rect 246304 336670 246356 336676
rect 246212 336592 246264 336598
rect 246212 336534 246264 336540
rect 246316 284986 246344 336670
rect 246592 328574 246620 338014
rect 247098 337770 247126 338028
rect 247236 338014 247480 338042
rect 247604 338014 247848 338042
rect 247972 338014 248216 338042
rect 248432 338014 248584 338042
rect 248708 338014 248952 338042
rect 249076 338014 249320 338042
rect 249444 338014 249688 338042
rect 249996 338014 250056 338042
rect 250180 338014 250424 338042
rect 250548 338014 250792 338042
rect 250916 338014 251160 338042
rect 251284 338014 251528 338042
rect 251652 338014 251896 338042
rect 252020 338014 252264 338042
rect 247098 337742 247172 337770
rect 246580 328568 246632 328574
rect 246580 328510 246632 328516
rect 246304 284980 246356 284986
rect 246304 284922 246356 284928
rect 246396 4820 246448 4826
rect 246396 4762 246448 4768
rect 245936 3936 245988 3942
rect 245936 3878 245988 3884
rect 246408 480 246436 4762
rect 247144 4010 247172 337742
rect 247236 336734 247264 338014
rect 247224 336728 247276 336734
rect 247224 336670 247276 336676
rect 247604 335354 247632 338014
rect 247328 335326 247632 335354
rect 247328 330562 247356 335326
rect 247236 330534 247356 330562
rect 247236 207670 247264 330534
rect 247972 316034 248000 338014
rect 248432 320822 248460 338014
rect 248708 330426 248736 338014
rect 248524 330398 248736 330426
rect 248420 320816 248472 320822
rect 248420 320758 248472 320764
rect 247328 316006 248000 316034
rect 247224 207664 247276 207670
rect 247224 207606 247276 207612
rect 247224 31068 247276 31074
rect 247224 31010 247276 31016
rect 247132 4004 247184 4010
rect 247132 3946 247184 3952
rect 247236 3482 247264 31010
rect 247328 4078 247356 316006
rect 248524 64190 248552 330398
rect 248604 320816 248656 320822
rect 248604 320758 248656 320764
rect 248616 224262 248644 320758
rect 249076 316034 249104 338014
rect 249444 331906 249472 338014
rect 249432 331900 249484 331906
rect 249432 331842 249484 331848
rect 249800 330540 249852 330546
rect 249800 330482 249852 330488
rect 248708 316006 249104 316034
rect 248604 224256 248656 224262
rect 248604 224198 248656 224204
rect 248512 64184 248564 64190
rect 248512 64126 248564 64132
rect 248512 22840 248564 22846
rect 248512 22782 248564 22788
rect 247316 4072 247368 4078
rect 247316 4014 247368 4020
rect 247236 3454 247632 3482
rect 247604 480 247632 3454
rect 240478 354 240590 480
rect 240336 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248524 354 248552 22782
rect 248708 4146 248736 316006
rect 249812 50386 249840 330482
rect 249892 330472 249944 330478
rect 249892 330414 249944 330420
rect 249904 220114 249932 330414
rect 249996 221474 250024 338014
rect 250180 330546 250208 338014
rect 250168 330540 250220 330546
rect 250168 330482 250220 330488
rect 250548 322250 250576 338014
rect 250916 330478 250944 338014
rect 251180 330540 251232 330546
rect 251180 330482 251232 330488
rect 250904 330472 250956 330478
rect 250904 330414 250956 330420
rect 250536 322244 250588 322250
rect 250536 322186 250588 322192
rect 249984 221468 250036 221474
rect 249984 221410 250036 221416
rect 249892 220108 249944 220114
rect 249892 220050 249944 220056
rect 249800 50380 249852 50386
rect 249800 50322 249852 50328
rect 251192 32434 251220 330482
rect 251284 61402 251312 338014
rect 251652 316034 251680 338014
rect 251824 336728 251876 336734
rect 251824 336670 251876 336676
rect 251376 316006 251680 316034
rect 251376 304298 251404 316006
rect 251364 304292 251416 304298
rect 251364 304234 251416 304240
rect 251836 217326 251864 336670
rect 252020 330546 252048 338014
rect 252618 337770 252646 338028
rect 252756 338014 253000 338042
rect 253124 338014 253368 338042
rect 253492 338014 253736 338042
rect 253952 338014 254104 338042
rect 254228 338014 254472 338042
rect 254596 338014 254840 338042
rect 254964 338014 255208 338042
rect 255516 338014 255576 338042
rect 255700 338014 255944 338042
rect 256068 338014 256312 338042
rect 256436 338014 256680 338042
rect 256896 338014 257048 338042
rect 257172 338014 257416 338042
rect 257540 338014 257784 338042
rect 258152 338014 258304 338042
rect 252618 337742 252692 337770
rect 252008 330540 252060 330546
rect 252008 330482 252060 330488
rect 251824 217320 251876 217326
rect 251824 217262 251876 217268
rect 252664 206310 252692 337742
rect 252756 330682 252784 338014
rect 253124 335354 253152 338014
rect 252848 335326 253152 335354
rect 252744 330676 252796 330682
rect 252744 330618 252796 330624
rect 252848 330562 252876 335326
rect 252756 330534 252876 330562
rect 252756 218754 252784 330534
rect 253492 316034 253520 338014
rect 253952 329118 253980 338014
rect 254228 336734 254256 338014
rect 254216 336728 254268 336734
rect 254216 336670 254268 336676
rect 254032 330540 254084 330546
rect 254032 330482 254084 330488
rect 253940 329112 253992 329118
rect 253940 329054 253992 329060
rect 252848 316006 253520 316034
rect 252744 218748 252796 218754
rect 252744 218690 252796 218696
rect 252652 206304 252704 206310
rect 252652 206246 252704 206252
rect 251272 61396 251324 61402
rect 251272 61338 251324 61344
rect 251272 50380 251324 50386
rect 251272 50322 251324 50328
rect 251180 32428 251232 32434
rect 251180 32370 251232 32376
rect 249800 18624 249852 18630
rect 249800 18566 249852 18572
rect 249812 16574 249840 18566
rect 249812 16546 250024 16574
rect 248696 4140 248748 4146
rect 248696 4082 248748 4088
rect 249996 480 250024 16546
rect 251284 3602 251312 50322
rect 251364 32428 251416 32434
rect 251364 32370 251416 32376
rect 251272 3596 251324 3602
rect 251272 3538 251324 3544
rect 251376 3482 251404 32370
rect 252848 22778 252876 316006
rect 254044 307086 254072 330482
rect 254596 316034 254624 338014
rect 254964 330546 254992 338014
rect 254952 330540 255004 330546
rect 254952 330482 255004 330488
rect 255412 330540 255464 330546
rect 255412 330482 255464 330488
rect 255320 330472 255372 330478
rect 255320 330414 255372 330420
rect 254228 316006 254624 316034
rect 254032 307080 254084 307086
rect 254032 307022 254084 307028
rect 254228 204950 254256 316006
rect 254216 204944 254268 204950
rect 254216 204886 254268 204892
rect 255332 51746 255360 330414
rect 255424 203590 255452 330482
rect 255516 215966 255544 338014
rect 255700 330546 255728 338014
rect 255688 330540 255740 330546
rect 255688 330482 255740 330488
rect 256068 316034 256096 338014
rect 256436 330478 256464 338014
rect 256700 330540 256752 330546
rect 256700 330482 256752 330488
rect 256424 330472 256476 330478
rect 256424 330414 256476 330420
rect 255608 316006 256096 316034
rect 255608 312594 255636 316006
rect 255596 312588 255648 312594
rect 255596 312530 255648 312536
rect 255504 215960 255556 215966
rect 255504 215902 255556 215908
rect 255412 203584 255464 203590
rect 255412 203526 255464 203532
rect 255320 51740 255372 51746
rect 255320 51682 255372 51688
rect 255412 51740 255464 51746
rect 255412 51682 255464 51688
rect 252836 22772 252888 22778
rect 252836 22714 252888 22720
rect 255424 16574 255452 51682
rect 255424 16546 255912 16574
rect 254216 11824 254268 11830
rect 254216 11766 254268 11772
rect 253480 9104 253532 9110
rect 253480 9046 253532 9052
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251192 3454 251404 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3538
rect 253492 480 253520 9046
rect 248758 354 248870 480
rect 248524 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 11766
rect 255884 480 255912 16546
rect 256712 8974 256740 330482
rect 256792 330472 256844 330478
rect 256792 330414 256844 330420
rect 256804 33794 256832 330414
rect 256896 202162 256924 338014
rect 257172 330546 257200 338014
rect 257160 330540 257212 330546
rect 257160 330482 257212 330488
rect 257540 330478 257568 338014
rect 258276 330562 258304 338014
rect 258460 338014 258520 338042
rect 258644 338014 258888 338042
rect 259012 338014 259164 338042
rect 259472 338014 259532 338042
rect 259656 338014 259900 338042
rect 260024 338014 260268 338042
rect 260392 338014 260636 338042
rect 258172 330540 258224 330546
rect 258276 330534 258396 330562
rect 258172 330482 258224 330488
rect 257528 330472 257580 330478
rect 257528 330414 257580 330420
rect 258080 330404 258132 330410
rect 258080 330346 258132 330352
rect 256884 202156 256936 202162
rect 256884 202098 256936 202104
rect 256792 33788 256844 33794
rect 256792 33730 256844 33736
rect 256792 21480 256844 21486
rect 256792 21422 256844 21428
rect 256700 8968 256752 8974
rect 256700 8910 256752 8916
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256804 354 256832 21422
rect 258092 9042 258120 330346
rect 258184 14482 258212 330482
rect 258264 330472 258316 330478
rect 258264 330414 258316 330420
rect 258276 200802 258304 330414
rect 258368 308446 258396 330534
rect 258460 330410 258488 338014
rect 258644 330546 258672 338014
rect 258632 330540 258684 330546
rect 258632 330482 258684 330488
rect 259012 330478 259040 338014
rect 259000 330472 259052 330478
rect 259000 330414 259052 330420
rect 258448 330404 258500 330410
rect 258448 330346 258500 330352
rect 258356 308440 258408 308446
rect 258356 308382 258408 308388
rect 258264 200796 258316 200802
rect 258264 200738 258316 200744
rect 258264 33788 258316 33794
rect 258264 33730 258316 33736
rect 258172 14476 258224 14482
rect 258172 14418 258224 14424
rect 258080 9036 258132 9042
rect 258080 8978 258132 8984
rect 258276 480 258304 33730
rect 259472 10334 259500 338014
rect 259552 327684 259604 327690
rect 259552 327626 259604 327632
rect 259564 10402 259592 327626
rect 259656 14550 259684 338014
rect 260024 316034 260052 338014
rect 260392 327690 260420 338014
rect 260990 337770 261018 338028
rect 261128 338014 261372 338042
rect 261496 338014 261740 338042
rect 261864 338014 262108 338042
rect 262416 338014 262476 338042
rect 262600 338014 262844 338042
rect 262968 338014 263212 338042
rect 263336 338014 263580 338042
rect 263704 338014 263948 338042
rect 264072 338014 264316 338042
rect 264440 338014 264684 338042
rect 264992 338014 265052 338042
rect 265176 338014 265420 338042
rect 265544 338014 265788 338042
rect 265912 338014 266156 338042
rect 266524 338014 266676 338042
rect 260990 337742 261064 337770
rect 260840 335980 260892 335986
rect 260840 335922 260892 335928
rect 260380 327684 260432 327690
rect 260380 327626 260432 327632
rect 259748 316006 260052 316034
rect 259748 289134 259776 316006
rect 259736 289128 259788 289134
rect 259736 289070 259788 289076
rect 260852 35222 260880 335922
rect 260932 330540 260984 330546
rect 260932 330482 260984 330488
rect 260944 213246 260972 330482
rect 261036 214606 261064 337742
rect 261128 335986 261156 338014
rect 261116 335980 261168 335986
rect 261116 335922 261168 335928
rect 261496 316034 261524 338014
rect 261864 330546 261892 338014
rect 261852 330540 261904 330546
rect 261852 330482 261904 330488
rect 262312 330540 262364 330546
rect 262312 330482 262364 330488
rect 262220 329316 262272 329322
rect 262220 329258 262272 329264
rect 261128 316006 261524 316034
rect 261128 276690 261156 316006
rect 261116 276684 261168 276690
rect 261116 276626 261168 276632
rect 261024 214600 261076 214606
rect 261024 214542 261076 214548
rect 260932 213240 260984 213246
rect 260932 213182 260984 213188
rect 260840 35216 260892 35222
rect 260840 35158 260892 35164
rect 259736 24200 259788 24206
rect 259736 24142 259788 24148
rect 259644 14544 259696 14550
rect 259644 14486 259696 14492
rect 259552 10396 259604 10402
rect 259552 10338 259604 10344
rect 259460 10328 259512 10334
rect 259460 10270 259512 10276
rect 259748 6914 259776 24142
rect 260656 15972 260708 15978
rect 260656 15914 260708 15920
rect 259472 6886 259776 6914
rect 259472 480 259500 6886
rect 260668 480 260696 15914
rect 262232 14618 262260 329258
rect 262324 198014 262352 330482
rect 262416 199442 262444 338014
rect 262600 316034 262628 338014
rect 262968 329322 262996 338014
rect 263336 330546 263364 338014
rect 263704 336682 263732 338014
rect 263612 336654 263732 336682
rect 263324 330540 263376 330546
rect 263324 330482 263376 330488
rect 262956 329316 263008 329322
rect 262956 329258 263008 329264
rect 262508 316006 262628 316034
rect 262508 278050 262536 316006
rect 262496 278044 262548 278050
rect 262496 277986 262548 277992
rect 262404 199436 262456 199442
rect 262404 199378 262456 199384
rect 262312 198008 262364 198014
rect 262312 197950 262364 197956
rect 262312 26988 262364 26994
rect 262312 26930 262364 26936
rect 262324 16574 262352 26930
rect 262324 16546 262536 16574
rect 262220 14612 262272 14618
rect 262220 14554 262272 14560
rect 261760 8968 261812 8974
rect 261760 8910 261812 8916
rect 261772 480 261800 8910
rect 257038 354 257150 480
rect 256804 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 263612 13122 263640 336654
rect 264072 335354 264100 338014
rect 264440 336682 264468 338014
rect 263704 335326 264100 335354
rect 264164 336654 264468 336682
rect 263704 14686 263732 335326
rect 264164 316034 264192 336654
rect 264992 336122 265020 338014
rect 264244 336116 264296 336122
rect 264244 336058 264296 336064
rect 264980 336116 265032 336122
rect 264980 336058 265032 336064
rect 263796 316006 264192 316034
rect 263796 196654 263824 316006
rect 264256 279478 264284 336058
rect 265176 335354 265204 338014
rect 265084 335326 265204 335354
rect 264244 279472 264296 279478
rect 264244 279414 264296 279420
rect 265084 211818 265112 335326
rect 265164 328024 265216 328030
rect 265164 327966 265216 327972
rect 265176 227050 265204 327966
rect 265544 316034 265572 338014
rect 265912 328030 265940 338014
rect 266544 330540 266596 330546
rect 266544 330482 266596 330488
rect 266452 330472 266504 330478
rect 266452 330414 266504 330420
rect 265900 328024 265952 328030
rect 265900 327966 265952 327972
rect 265268 316006 265572 316034
rect 265164 227044 265216 227050
rect 265164 226986 265216 226992
rect 265072 211812 265124 211818
rect 265072 211754 265124 211760
rect 263784 196648 263836 196654
rect 263784 196590 263836 196596
rect 265268 62830 265296 316006
rect 266464 210458 266492 330414
rect 266556 225622 266584 330482
rect 266544 225616 266596 225622
rect 266544 225558 266596 225564
rect 266452 210452 266504 210458
rect 266452 210394 266504 210400
rect 265256 62824 265308 62830
rect 265256 62766 265308 62772
rect 266648 60042 266676 338014
rect 266740 338014 266892 338042
rect 267016 338014 267260 338042
rect 267384 338014 267628 338042
rect 267936 338014 267996 338042
rect 268120 338014 268364 338042
rect 268488 338014 268732 338042
rect 268856 338014 269100 338042
rect 269224 338014 269468 338042
rect 269592 338014 269836 338042
rect 269960 338014 270204 338042
rect 266740 336054 266768 338014
rect 266728 336048 266780 336054
rect 266728 335990 266780 335996
rect 267016 330546 267044 338014
rect 267004 330540 267056 330546
rect 267004 330482 267056 330488
rect 267384 330478 267412 338014
rect 267832 330540 267884 330546
rect 267832 330482 267884 330488
rect 267372 330472 267424 330478
rect 267372 330414 267424 330420
rect 266636 60036 266688 60042
rect 266636 59978 266688 59984
rect 263784 22772 263836 22778
rect 263784 22714 263836 22720
rect 263796 16574 263824 22714
rect 263796 16546 264192 16574
rect 263692 14680 263744 14686
rect 263692 14622 263744 14628
rect 263600 13116 263652 13122
rect 263600 13058 263652 13064
rect 264164 480 264192 16546
rect 267844 14754 267872 330482
rect 267936 195294 267964 338014
rect 267924 195288 267976 195294
rect 267924 195230 267976 195236
rect 267924 35216 267976 35222
rect 267924 35158 267976 35164
rect 267832 14748 267884 14754
rect 267832 14690 267884 14696
rect 267740 14476 267792 14482
rect 267740 14418 267792 14424
rect 264980 10328 265032 10334
rect 264980 10270 265032 10276
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 10270
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 266556 480 266584 3470
rect 267752 480 267780 14418
rect 267936 6914 267964 35158
rect 268120 13190 268148 338014
rect 268488 330546 268516 338014
rect 268856 336190 268884 338014
rect 268844 336184 268896 336190
rect 268844 336126 268896 336132
rect 268476 330540 268528 330546
rect 268476 330482 268528 330488
rect 269120 330540 269172 330546
rect 269120 330482 269172 330488
rect 268108 13184 268160 13190
rect 268108 13126 268160 13132
rect 267936 6886 268424 6914
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 6886
rect 269132 3398 269160 330482
rect 269224 13258 269252 338014
rect 269592 316034 269620 338014
rect 269764 336728 269816 336734
rect 269764 336670 269816 336676
rect 269776 327758 269804 336670
rect 269960 330546 269988 338014
rect 270558 337822 270586 338028
rect 270546 337816 270598 337822
rect 270546 337758 270598 337764
rect 269948 330540 270000 330546
rect 269948 330482 270000 330488
rect 270592 330540 270644 330546
rect 270592 330482 270644 330488
rect 269764 327752 269816 327758
rect 269764 327694 269816 327700
rect 269316 316006 269620 316034
rect 269316 14822 269344 316006
rect 269304 14816 269356 14822
rect 269304 14758 269356 14764
rect 270604 13394 270632 330482
rect 270696 15910 270724 338150
rect 271064 338014 271216 338042
rect 271340 338014 271584 338042
rect 271952 338014 272104 338042
rect 270776 337816 270828 337822
rect 270776 337758 270828 337764
rect 270684 15904 270736 15910
rect 270684 15846 270736 15852
rect 270592 13388 270644 13394
rect 270592 13330 270644 13336
rect 270788 13326 270816 337758
rect 271064 336258 271092 338014
rect 271052 336252 271104 336258
rect 271052 336194 271104 336200
rect 271144 335844 271196 335850
rect 271144 335786 271196 335792
rect 271156 280838 271184 335786
rect 271340 330546 271368 338014
rect 271328 330540 271380 330546
rect 271328 330482 271380 330488
rect 271972 330540 272024 330546
rect 271972 330482 272024 330488
rect 271984 311166 272012 330482
rect 272076 313954 272104 338014
rect 272168 338014 272320 338042
rect 272444 338014 272688 338042
rect 272812 338014 273056 338042
rect 272064 313948 272116 313954
rect 272064 313890 272116 313896
rect 271972 311160 272024 311166
rect 271972 311102 272024 311108
rect 271144 280832 271196 280838
rect 271144 280774 271196 280780
rect 270776 13320 270828 13326
rect 270776 13262 270828 13268
rect 269212 13252 269264 13258
rect 269212 13194 269264 13200
rect 270776 13116 270828 13122
rect 270776 13058 270828 13064
rect 269120 3392 269172 3398
rect 269120 3334 269172 3340
rect 270040 3188 270092 3194
rect 270040 3130 270092 3136
rect 270052 480 270080 3130
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 13058
rect 272168 3330 272196 338014
rect 272444 335850 272472 338014
rect 272432 335844 272484 335850
rect 272432 335786 272484 335792
rect 272812 330546 272840 338014
rect 273410 337770 273438 338028
rect 273548 338014 273792 338042
rect 273916 338014 274160 338042
rect 274284 338014 274528 338042
rect 274836 338014 274896 338042
rect 275020 338014 275264 338042
rect 275388 338014 275632 338042
rect 275756 338014 276000 338042
rect 276124 338014 276368 338042
rect 276492 338014 276736 338042
rect 276860 338014 277104 338042
rect 277472 338014 277624 338042
rect 273410 337742 273484 337770
rect 272800 330540 272852 330546
rect 272800 330482 272852 330488
rect 273352 322108 273404 322114
rect 273352 322050 273404 322056
rect 273364 24138 273392 322050
rect 273352 24132 273404 24138
rect 273352 24074 273404 24080
rect 272432 7744 272484 7750
rect 272432 7686 272484 7692
rect 272156 3324 272208 3330
rect 272156 3266 272208 3272
rect 272444 480 272472 7686
rect 273456 3262 273484 337742
rect 273548 336734 273576 338014
rect 273536 336728 273588 336734
rect 273536 336670 273588 336676
rect 273916 322114 273944 338014
rect 274284 336394 274312 338014
rect 274272 336388 274324 336394
rect 274272 336330 274324 336336
rect 274640 326392 274692 326398
rect 274640 326334 274692 326340
rect 273904 322108 273956 322114
rect 273904 322050 273956 322056
rect 274652 273970 274680 326334
rect 274836 323678 274864 338014
rect 275020 326398 275048 338014
rect 275388 331214 275416 338014
rect 275112 331186 275416 331214
rect 275008 326392 275060 326398
rect 275008 326334 275060 326340
rect 274824 323672 274876 323678
rect 274824 323614 274876 323620
rect 275112 323490 275140 331186
rect 274744 323462 275140 323490
rect 274640 273964 274692 273970
rect 274640 273906 274692 273912
rect 274744 233918 274772 323462
rect 275756 321554 275784 338014
rect 276020 326392 276072 326398
rect 276020 326334 276072 326340
rect 274836 321526 275784 321554
rect 274836 308514 274864 321526
rect 274824 308508 274876 308514
rect 274824 308450 274876 308456
rect 274824 274100 274876 274106
rect 274824 274042 274876 274048
rect 274732 233912 274784 233918
rect 274732 233854 274784 233860
rect 273628 3596 273680 3602
rect 273628 3538 273680 3544
rect 273444 3256 273496 3262
rect 273444 3198 273496 3204
rect 273640 480 273668 3538
rect 274836 480 274864 274042
rect 276032 54534 276060 326334
rect 276124 250510 276152 338014
rect 276492 326398 276520 338014
rect 276860 336682 276888 338014
rect 276584 336654 276888 336682
rect 276480 326392 276532 326398
rect 276480 326334 276532 326340
rect 276584 316034 276612 336654
rect 276664 336252 276716 336258
rect 276664 336194 276716 336200
rect 276216 316006 276612 316034
rect 276216 309806 276244 316006
rect 276204 309800 276256 309806
rect 276204 309742 276256 309748
rect 276676 287706 276704 336194
rect 276756 336048 276808 336054
rect 276756 335990 276808 335996
rect 276768 324970 276796 335990
rect 277492 326392 277544 326398
rect 277492 326334 277544 326340
rect 276756 324964 276808 324970
rect 276756 324906 276808 324912
rect 276664 287700 276716 287706
rect 276664 287642 276716 287648
rect 276204 250640 276256 250646
rect 276204 250582 276256 250588
rect 276112 250504 276164 250510
rect 276112 250446 276164 250452
rect 276020 54528 276072 54534
rect 276020 54470 276072 54476
rect 276216 6914 276244 250582
rect 277504 247722 277532 326334
rect 277596 290494 277624 338014
rect 277688 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278576 338042
rect 278884 338014 278944 338042
rect 279068 338014 279312 338042
rect 279436 338014 279680 338042
rect 279804 338014 280048 338042
rect 277584 290488 277636 290494
rect 277584 290430 277636 290436
rect 277492 247716 277544 247722
rect 277492 247658 277544 247664
rect 277688 36582 277716 338014
rect 277964 336258 277992 338014
rect 277952 336252 278004 336258
rect 277952 336194 278004 336200
rect 278332 326398 278360 338014
rect 278320 326392 278372 326398
rect 278320 326334 278372 326340
rect 278780 326324 278832 326330
rect 278780 326266 278832 326272
rect 277676 36576 277728 36582
rect 277676 36518 277728 36524
rect 278792 21418 278820 326266
rect 278884 228410 278912 338014
rect 278964 326392 279016 326398
rect 278964 326334 279016 326340
rect 278976 246362 279004 326334
rect 279068 300150 279096 338014
rect 279436 326398 279464 338014
rect 279424 326392 279476 326398
rect 279424 326334 279476 326340
rect 279804 326330 279832 338014
rect 280402 337770 280430 338028
rect 280540 338014 280784 338042
rect 280908 338014 281152 338042
rect 281276 338014 281520 338042
rect 281644 338014 281888 338042
rect 282012 338014 282256 338042
rect 282380 338014 282624 338042
rect 282992 338014 283144 338042
rect 280402 337742 280476 337770
rect 280448 331226 280476 337742
rect 280436 331220 280488 331226
rect 280436 331162 280488 331168
rect 280540 326618 280568 338014
rect 280620 331220 280672 331226
rect 280620 331162 280672 331168
rect 280264 326590 280568 326618
rect 279792 326324 279844 326330
rect 279792 326266 279844 326272
rect 280160 326324 280212 326330
rect 280160 326266 280212 326272
rect 279056 300144 279108 300150
rect 279056 300086 279108 300092
rect 278964 246356 279016 246362
rect 278964 246298 279016 246304
rect 278872 228404 278924 228410
rect 278872 228346 278924 228352
rect 280172 53106 280200 326266
rect 280264 244934 280292 326590
rect 280344 326392 280396 326398
rect 280344 326334 280396 326340
rect 280356 272542 280384 326334
rect 280632 316034 280660 331162
rect 280908 326330 280936 338014
rect 281276 326398 281304 338014
rect 281264 326392 281316 326398
rect 281264 326334 281316 326340
rect 281540 326392 281592 326398
rect 281540 326334 281592 326340
rect 280896 326324 280948 326330
rect 280896 326266 280948 326272
rect 280448 316006 280660 316034
rect 280448 301510 280476 316006
rect 280436 301504 280488 301510
rect 280436 301446 280488 301452
rect 280344 272536 280396 272542
rect 280344 272478 280396 272484
rect 280252 244928 280304 244934
rect 280252 244870 280304 244876
rect 281552 55894 281580 326334
rect 281644 243574 281672 338014
rect 282012 326398 282040 338014
rect 282000 326392 282052 326398
rect 282000 326334 282052 326340
rect 282380 316034 282408 338014
rect 282828 336728 282880 336734
rect 282828 336670 282880 336676
rect 282840 329186 282868 336670
rect 283116 335354 283144 338014
rect 283254 337770 283282 338028
rect 283392 338014 283636 338042
rect 283760 338014 284004 338042
rect 283254 337742 283328 337770
rect 283116 335326 283236 335354
rect 283208 330818 283236 335326
rect 283196 330812 283248 330818
rect 283196 330754 283248 330760
rect 283300 330698 283328 337742
rect 282932 330670 283328 330698
rect 282828 329180 282880 329186
rect 282828 329122 282880 329128
rect 281736 316006 282408 316034
rect 281736 271182 281764 316006
rect 281724 271176 281776 271182
rect 281724 271118 281776 271124
rect 281632 243568 281684 243574
rect 281632 243510 281684 243516
rect 282932 57254 282960 330670
rect 283392 330562 283420 338014
rect 283472 330812 283524 330818
rect 283472 330754 283524 330760
rect 283116 330534 283420 330562
rect 283012 329180 283064 329186
rect 283012 329122 283064 329128
rect 283024 242214 283052 329122
rect 283116 289202 283144 330534
rect 283484 330426 283512 330754
rect 283208 330398 283512 330426
rect 283208 291854 283236 330398
rect 283760 329186 283788 338014
rect 284358 337770 284386 338028
rect 284496 338014 284740 338042
rect 284864 338014 285108 338042
rect 285232 338014 285476 338042
rect 285692 338014 285844 338042
rect 285968 338014 286212 338042
rect 286336 338014 286580 338042
rect 286704 338014 286948 338042
rect 287256 338014 287316 338042
rect 287440 338014 287684 338042
rect 287808 338014 288052 338042
rect 288176 338014 288420 338042
rect 288544 338014 288788 338042
rect 288912 338014 289156 338042
rect 289280 338014 289524 338042
rect 284358 337742 284432 337770
rect 283748 329180 283800 329186
rect 283748 329122 283800 329128
rect 283196 291848 283248 291854
rect 283196 291790 283248 291796
rect 283104 289196 283156 289202
rect 283104 289138 283156 289144
rect 283012 242208 283064 242214
rect 283012 242150 283064 242156
rect 284404 58682 284432 337742
rect 284496 336054 284524 338014
rect 284484 336048 284536 336054
rect 284484 335990 284536 335996
rect 284864 335354 284892 338014
rect 284496 335326 284892 335354
rect 284496 269822 284524 335326
rect 285232 316034 285260 338014
rect 285692 336734 285720 338014
rect 285680 336728 285732 336734
rect 285680 336670 285732 336676
rect 285772 330540 285824 330546
rect 285772 330482 285824 330488
rect 284588 316006 285260 316034
rect 284484 269816 284536 269822
rect 284484 269758 284536 269764
rect 284392 58676 284444 58682
rect 284392 58618 284444 58624
rect 282920 57248 282972 57254
rect 282920 57190 282972 57196
rect 281540 55888 281592 55894
rect 281540 55830 281592 55836
rect 280160 53100 280212 53106
rect 280160 53042 280212 53048
rect 282920 36576 282972 36582
rect 282920 36518 282972 36524
rect 281540 24132 281592 24138
rect 281540 24074 281592 24080
rect 278780 21412 278832 21418
rect 278780 21354 278832 21360
rect 279056 15904 279108 15910
rect 279056 15846 279108 15852
rect 276032 6886 276244 6914
rect 276032 480 276060 6886
rect 278320 4888 278372 4894
rect 278320 4830 278372 4836
rect 277122 3360 277178 3369
rect 277122 3295 277178 3304
rect 277136 480 277164 3295
rect 278332 480 278360 4830
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 15846
rect 280712 3664 280764 3670
rect 280712 3606 280764 3612
rect 280724 480 280752 3606
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 24074
rect 282932 16574 282960 36518
rect 284588 25634 284616 316006
rect 285680 284980 285732 284986
rect 285680 284922 285732 284928
rect 284576 25628 284628 25634
rect 284576 25570 284628 25576
rect 284392 25560 284444 25566
rect 284392 25502 284444 25508
rect 284404 16574 284432 25502
rect 285692 16574 285720 284922
rect 285784 239426 285812 330482
rect 285968 316034 285996 338014
rect 286232 336048 286284 336054
rect 286232 335990 286284 335996
rect 286244 325694 286272 335990
rect 286336 330546 286364 338014
rect 286416 335776 286468 335782
rect 286416 335718 286468 335724
rect 286324 330540 286376 330546
rect 286324 330482 286376 330488
rect 286244 325666 286364 325694
rect 285876 316006 285996 316034
rect 285876 268394 285904 316006
rect 286336 285054 286364 325666
rect 286428 312662 286456 335718
rect 286704 330614 286732 338014
rect 286692 330608 286744 330614
rect 286692 330550 286744 330556
rect 287152 330540 287204 330546
rect 287152 330482 287204 330488
rect 286416 312656 286468 312662
rect 286416 312598 286468 312604
rect 286324 285048 286376 285054
rect 286324 284990 286376 284996
rect 285864 268388 285916 268394
rect 285864 268330 285916 268336
rect 287164 264246 287192 330482
rect 287256 265674 287284 338014
rect 287440 316034 287468 338014
rect 287704 336728 287756 336734
rect 287704 336670 287756 336676
rect 287348 316006 287468 316034
rect 287244 265668 287296 265674
rect 287244 265610 287296 265616
rect 287152 264240 287204 264246
rect 287152 264182 287204 264188
rect 285772 239420 285824 239426
rect 285772 239362 285824 239368
rect 287348 37942 287376 316006
rect 287716 303006 287744 336670
rect 287808 335782 287836 338014
rect 287796 335776 287848 335782
rect 287796 335718 287848 335724
rect 288176 330546 288204 338014
rect 288164 330540 288216 330546
rect 288164 330482 288216 330488
rect 287704 303000 287756 303006
rect 287704 302942 287756 302948
rect 287336 37936 287388 37942
rect 287336 37878 287388 37884
rect 282932 16546 283144 16574
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 283116 480 283144 16546
rect 284300 3732 284352 3738
rect 284300 3674 284352 3680
rect 284312 480 284340 3674
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 288544 10470 288572 338014
rect 288912 331974 288940 338014
rect 289280 336682 289308 338014
rect 289878 337770 289906 338028
rect 290016 338014 290260 338042
rect 290384 338014 290628 338042
rect 290752 338014 290996 338042
rect 291212 338014 291364 338042
rect 291488 338014 291732 338042
rect 291856 338014 292100 338042
rect 292224 338014 292468 338042
rect 292592 338014 292836 338042
rect 292960 338014 293204 338042
rect 293328 338014 293572 338042
rect 293696 338014 293940 338042
rect 294064 338014 294308 338042
rect 294432 338014 294676 338042
rect 294800 338014 295044 338042
rect 295168 338014 295320 338042
rect 295536 338014 295688 338042
rect 295812 338014 296056 338042
rect 296180 338014 296424 338042
rect 296732 338014 296792 338042
rect 296916 338014 297160 338042
rect 297284 338014 297528 338042
rect 297652 338014 297896 338042
rect 298204 338014 298264 338042
rect 298388 338014 298632 338042
rect 298756 338014 299000 338042
rect 299124 338014 299368 338042
rect 299676 338014 299736 338042
rect 299860 338014 300104 338042
rect 300228 338014 300472 338042
rect 300596 338014 300840 338042
rect 300964 338014 301208 338042
rect 301332 338014 301576 338042
rect 301700 338014 301944 338042
rect 302252 338014 302312 338042
rect 302436 338014 302680 338042
rect 302804 338014 303048 338042
rect 303172 338014 303416 338042
rect 303724 338014 303784 338042
rect 303908 338014 304152 338042
rect 304276 338014 304520 338042
rect 304644 338014 304888 338042
rect 289878 337742 289952 337770
rect 289004 336654 289308 336682
rect 288900 331968 288952 331974
rect 288900 331910 288952 331916
rect 289004 316034 289032 336654
rect 289084 336116 289136 336122
rect 289084 336058 289136 336064
rect 288728 316006 289032 316034
rect 288532 10464 288584 10470
rect 288532 10406 288584 10412
rect 288728 7614 288756 316006
rect 288992 10396 289044 10402
rect 288992 10338 289044 10344
rect 288716 7608 288768 7614
rect 288716 7550 288768 7556
rect 287796 3800 287848 3806
rect 287796 3742 287848 3748
rect 287808 480 287836 3742
rect 289004 480 289032 10338
rect 289096 4826 289124 336058
rect 289176 335572 289228 335578
rect 289176 335514 289228 335520
rect 289188 286414 289216 335514
rect 289924 325038 289952 337742
rect 290016 335578 290044 338014
rect 290384 336734 290412 338014
rect 290372 336728 290424 336734
rect 290372 336670 290424 336676
rect 290004 335572 290056 335578
rect 290004 335514 290056 335520
rect 289912 325032 289964 325038
rect 289912 324974 289964 324980
rect 290752 316034 290780 338014
rect 291212 336054 291240 338014
rect 291200 336048 291252 336054
rect 291200 335990 291252 335996
rect 291488 335354 291516 338014
rect 291856 336682 291884 338014
rect 290016 316006 290780 316034
rect 291304 335326 291516 335354
rect 291672 336654 291884 336682
rect 291936 336660 291988 336666
rect 289176 286408 289228 286414
rect 289176 286350 289228 286356
rect 290016 238066 290044 316006
rect 291304 262886 291332 335326
rect 291384 330540 291436 330546
rect 291384 330482 291436 330488
rect 291396 283694 291424 330482
rect 291672 316034 291700 336654
rect 291936 336602 291988 336608
rect 291844 336048 291896 336054
rect 291844 335990 291896 335996
rect 291488 316006 291700 316034
rect 291384 283688 291436 283694
rect 291384 283630 291436 283636
rect 291292 262880 291344 262886
rect 291292 262822 291344 262828
rect 290004 238060 290056 238066
rect 290004 238002 290056 238008
rect 291488 39370 291516 316006
rect 291476 39364 291528 39370
rect 291476 39306 291528 39312
rect 289820 18692 289872 18698
rect 289820 18634 289872 18640
rect 289084 4820 289136 4826
rect 289084 4762 289136 4768
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 18634
rect 291856 15978 291884 335990
rect 291948 322318 291976 336602
rect 292224 330546 292252 338014
rect 292212 330540 292264 330546
rect 292212 330482 292264 330488
rect 292592 324902 292620 338014
rect 292960 335354 292988 338014
rect 293224 336728 293276 336734
rect 293224 336670 293276 336676
rect 292868 335326 292988 335354
rect 292868 330426 292896 335326
rect 292684 330398 292896 330426
rect 292580 324896 292632 324902
rect 292580 324838 292632 324844
rect 291936 322312 291988 322318
rect 291936 322254 291988 322260
rect 292580 261588 292632 261594
rect 292580 261530 292632 261536
rect 292592 16574 292620 261530
rect 292684 236706 292712 330398
rect 293236 326466 293264 336670
rect 293328 336666 293356 338014
rect 293316 336660 293368 336666
rect 293316 336602 293368 336608
rect 293224 326460 293276 326466
rect 293224 326402 293276 326408
rect 292764 324896 292816 324902
rect 292764 324838 292816 324844
rect 292776 261526 292804 324838
rect 293696 316034 293724 338014
rect 292868 316006 293724 316034
rect 292764 261520 292816 261526
rect 292764 261462 292816 261468
rect 292868 260166 292896 316006
rect 292856 260160 292908 260166
rect 292856 260102 292908 260108
rect 292672 236700 292724 236706
rect 292672 236642 292724 236648
rect 294064 235278 294092 338014
rect 294432 336802 294460 338014
rect 294420 336796 294472 336802
rect 294420 336738 294472 336744
rect 294800 336682 294828 338014
rect 294156 336654 294828 336682
rect 294156 258806 294184 336654
rect 294604 336592 294656 336598
rect 294604 336534 294656 336540
rect 294236 330540 294288 330546
rect 294236 330482 294288 330488
rect 294144 258800 294196 258806
rect 294144 258742 294196 258748
rect 294052 235272 294104 235278
rect 294052 235214 294104 235220
rect 294248 40730 294276 330482
rect 294616 307154 294644 336534
rect 295168 330546 295196 338014
rect 295156 330540 295208 330546
rect 295156 330482 295208 330488
rect 295340 330540 295392 330546
rect 295340 330482 295392 330488
rect 294604 307148 294656 307154
rect 294604 307090 294656 307096
rect 294236 40724 294288 40730
rect 294236 40666 294288 40672
rect 292592 16546 293264 16574
rect 291844 15972 291896 15978
rect 291844 15914 291896 15920
rect 292580 4820 292632 4826
rect 292580 4762 292632 4768
rect 291384 3868 291436 3874
rect 291384 3810 291436 3816
rect 291396 480 291424 3810
rect 292592 480 292620 4762
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 295352 7682 295380 330482
rect 295432 328772 295484 328778
rect 295432 328714 295484 328720
rect 295444 42090 295472 328714
rect 295536 282266 295564 338014
rect 295812 330546 295840 338014
rect 295984 335368 296036 335374
rect 295984 335310 296036 335316
rect 295800 330540 295852 330546
rect 295800 330482 295852 330488
rect 295524 282260 295576 282266
rect 295524 282202 295576 282208
rect 295996 280906 296024 335310
rect 296180 328778 296208 338014
rect 296732 335374 296760 338014
rect 296720 335368 296772 335374
rect 296916 335354 296944 338014
rect 297284 335354 297312 338014
rect 297364 336184 297416 336190
rect 297364 336126 297416 336132
rect 296720 335310 296772 335316
rect 296824 335326 296944 335354
rect 297008 335326 297312 335354
rect 296824 330698 296852 335326
rect 296732 330670 296852 330698
rect 296168 328772 296220 328778
rect 296168 328714 296220 328720
rect 296732 327826 296760 330670
rect 297008 330528 297036 335326
rect 296824 330500 297036 330528
rect 296720 327820 296772 327826
rect 296720 327762 296772 327768
rect 295984 280900 296036 280906
rect 295984 280842 296036 280848
rect 296720 279676 296772 279682
rect 296720 279618 296772 279624
rect 295432 42084 295484 42090
rect 295432 42026 295484 42032
rect 296732 16574 296760 279618
rect 296824 232558 296852 330500
rect 296996 330404 297048 330410
rect 296996 330346 297048 330352
rect 297008 279546 297036 330346
rect 296996 279540 297048 279546
rect 296996 279482 297048 279488
rect 296812 232552 296864 232558
rect 296812 232494 296864 232500
rect 297376 18630 297404 336126
rect 297456 335708 297508 335714
rect 297456 335650 297508 335656
rect 297468 304366 297496 335650
rect 297652 330410 297680 338014
rect 297640 330404 297692 330410
rect 297640 330346 297692 330352
rect 297456 304360 297508 304366
rect 297456 304302 297508 304308
rect 298204 257446 298232 338014
rect 298388 335354 298416 338014
rect 298756 336666 298784 338014
rect 298744 336660 298796 336666
rect 298744 336602 298796 336608
rect 298744 336524 298796 336530
rect 298744 336466 298796 336472
rect 298296 335326 298416 335354
rect 298296 319462 298324 335326
rect 298376 330540 298428 330546
rect 298376 330482 298428 330488
rect 298284 319456 298336 319462
rect 298284 319398 298336 319404
rect 298192 257440 298244 257446
rect 298192 257382 298244 257388
rect 298388 256086 298416 330482
rect 298376 256080 298428 256086
rect 298376 256022 298428 256028
rect 298756 26926 298784 336466
rect 299124 330546 299152 338014
rect 299112 330540 299164 330546
rect 299112 330482 299164 330488
rect 299572 330540 299624 330546
rect 299572 330482 299624 330488
rect 299480 254788 299532 254794
rect 299480 254730 299532 254736
rect 298744 26920 298796 26926
rect 298744 26862 298796 26868
rect 297364 18624 297416 18630
rect 297364 18566 297416 18572
rect 296732 16546 297312 16574
rect 295340 7676 295392 7682
rect 295340 7618 295392 7624
rect 296076 4956 296128 4962
rect 296076 4898 296128 4904
rect 294880 3936 294932 3942
rect 294880 3878 294932 3884
rect 294892 480 294920 3878
rect 296088 480 296116 4898
rect 297284 480 297312 16546
rect 298468 4004 298520 4010
rect 298468 3946 298520 3952
rect 298480 480 298508 3946
rect 299492 3466 299520 254730
rect 299584 229770 299612 330482
rect 299676 231130 299704 338014
rect 299860 335714 299888 338014
rect 299848 335708 299900 335714
rect 299848 335650 299900 335656
rect 300228 316034 300256 338014
rect 300596 330546 300624 338014
rect 300768 336728 300820 336734
rect 300768 336670 300820 336676
rect 300780 334694 300808 336670
rect 300768 334688 300820 334694
rect 300768 334630 300820 334636
rect 300584 330540 300636 330546
rect 300584 330482 300636 330488
rect 300860 330540 300912 330546
rect 300860 330482 300912 330488
rect 299768 316006 300256 316034
rect 299768 254658 299796 316006
rect 299756 254652 299808 254658
rect 299756 254594 299808 254600
rect 299664 231124 299716 231130
rect 299664 231066 299716 231072
rect 299572 229764 299624 229770
rect 299572 229706 299624 229712
rect 300872 43450 300900 330482
rect 300964 278118 300992 338014
rect 301332 320890 301360 338014
rect 301504 335436 301556 335442
rect 301504 335378 301556 335384
rect 301320 320884 301372 320890
rect 301320 320826 301372 320832
rect 300952 278112 301004 278118
rect 300952 278054 301004 278060
rect 300860 43444 300912 43450
rect 300860 43386 300912 43392
rect 301516 11762 301544 335378
rect 301700 330546 301728 338014
rect 302252 336326 302280 338014
rect 302436 336530 302464 338014
rect 302424 336524 302476 336530
rect 302424 336466 302476 336472
rect 302240 336320 302292 336326
rect 302240 336262 302292 336268
rect 302804 335354 302832 338014
rect 302976 336524 303028 336530
rect 302976 336466 303028 336472
rect 302884 336252 302936 336258
rect 302884 336194 302936 336200
rect 302344 335326 302832 335354
rect 301688 330540 301740 330546
rect 301688 330482 301740 330488
rect 302344 318102 302372 335326
rect 302424 323332 302476 323338
rect 302424 323274 302476 323280
rect 302332 318096 302384 318102
rect 302332 318038 302384 318044
rect 302436 276758 302464 323274
rect 302424 276752 302476 276758
rect 302424 276694 302476 276700
rect 301504 11756 301556 11762
rect 301504 11698 301556 11704
rect 302896 10334 302924 336194
rect 302988 17338 303016 336466
rect 303172 323338 303200 338014
rect 303528 335640 303580 335646
rect 303528 335582 303580 335588
rect 303540 333266 303568 335582
rect 303528 333260 303580 333266
rect 303528 333202 303580 333208
rect 303160 323332 303212 323338
rect 303160 323274 303212 323280
rect 303724 267034 303752 338014
rect 303908 335354 303936 338014
rect 304276 336818 304304 338014
rect 304092 336790 304304 336818
rect 304092 336734 304120 336790
rect 304080 336728 304132 336734
rect 304644 336682 304672 338014
rect 305242 337770 305270 338028
rect 305380 338014 305624 338042
rect 305748 338014 305992 338042
rect 306116 338014 306360 338042
rect 306484 338014 306728 338042
rect 306852 338014 307096 338042
rect 307220 338014 307372 338042
rect 307496 338014 307740 338042
rect 307864 338014 308108 338042
rect 308232 338014 308476 338042
rect 308600 338014 308844 338042
rect 305242 337742 305316 337770
rect 304080 336670 304132 336676
rect 303816 335326 303936 335354
rect 304184 336654 304672 336682
rect 303816 316742 303844 335326
rect 303804 316736 303856 316742
rect 303804 316678 303856 316684
rect 304184 316034 304212 336654
rect 304264 335368 304316 335374
rect 304264 335310 304316 335316
rect 303908 316006 304212 316034
rect 303712 267028 303764 267034
rect 303712 266970 303764 266976
rect 303620 253428 303672 253434
rect 303620 253370 303672 253376
rect 302976 17332 303028 17338
rect 302976 17274 303028 17280
rect 303632 16574 303660 253370
rect 303908 253298 303936 316006
rect 303896 253292 303948 253298
rect 303896 253234 303948 253240
rect 303632 16546 303936 16574
rect 302884 10328 302936 10334
rect 302884 10270 302936 10276
rect 303160 5092 303212 5098
rect 303160 5034 303212 5040
rect 299664 5024 299716 5030
rect 299664 4966 299716 4972
rect 299480 3460 299532 3466
rect 299480 3402 299532 3408
rect 299676 480 299704 4966
rect 301964 4072 302016 4078
rect 301964 4014 302016 4020
rect 300768 3460 300820 3466
rect 300768 3402 300820 3408
rect 300780 480 300808 3402
rect 301976 480 302004 4014
rect 303172 480 303200 5034
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304276 6254 304304 335310
rect 305288 328454 305316 337742
rect 305196 328426 305316 328454
rect 305000 326392 305052 326398
rect 305000 326334 305052 326340
rect 305012 44878 305040 326334
rect 305196 323762 305224 328426
rect 305196 323734 305316 323762
rect 305184 323604 305236 323610
rect 305184 323546 305236 323552
rect 305092 322516 305144 322522
rect 305092 322458 305144 322464
rect 305104 251938 305132 322458
rect 305196 275398 305224 323546
rect 305288 315314 305316 323734
rect 305380 323610 305408 338014
rect 305644 335980 305696 335986
rect 305644 335922 305696 335928
rect 305368 323604 305420 323610
rect 305368 323546 305420 323552
rect 305276 315308 305328 315314
rect 305276 315250 305328 315256
rect 305184 275392 305236 275398
rect 305184 275334 305236 275340
rect 305092 251932 305144 251938
rect 305092 251874 305144 251880
rect 305656 46238 305684 335922
rect 305748 322522 305776 338014
rect 306116 326398 306144 338014
rect 306484 335646 306512 338014
rect 306472 335640 306524 335646
rect 306472 335582 306524 335588
rect 306852 335354 306880 338014
rect 307024 336728 307076 336734
rect 307024 336670 307076 336676
rect 306484 335326 306880 335354
rect 306104 326392 306156 326398
rect 306104 326334 306156 326340
rect 305736 322516 305788 322522
rect 305736 322458 305788 322464
rect 306484 249150 306512 335326
rect 306564 326392 306616 326398
rect 306564 326334 306616 326340
rect 306472 249144 306524 249150
rect 306472 249086 306524 249092
rect 305644 46232 305696 46238
rect 305644 46174 305696 46180
rect 305000 44872 305052 44878
rect 305000 44814 305052 44820
rect 306576 6322 306604 326334
rect 307036 11830 307064 336670
rect 307116 336660 307168 336666
rect 307116 336602 307168 336608
rect 307128 24206 307156 336602
rect 307220 335986 307248 338014
rect 307208 335980 307260 335986
rect 307208 335922 307260 335928
rect 307496 326398 307524 338014
rect 307864 335374 307892 338014
rect 307852 335368 307904 335374
rect 307852 335310 307904 335316
rect 307484 326392 307536 326398
rect 307484 326334 307536 326340
rect 308232 316034 308260 338014
rect 308600 335442 308628 338014
rect 309198 337770 309226 338028
rect 309428 338014 309580 338042
rect 309704 338014 309948 338042
rect 310072 338014 310316 338042
rect 309198 337742 309272 337770
rect 308588 335436 308640 335442
rect 308588 335378 308640 335384
rect 307864 316006 308260 316034
rect 307864 47598 307892 316006
rect 307852 47592 307904 47598
rect 307852 47534 307904 47540
rect 309244 28286 309272 337742
rect 309324 326392 309376 326398
rect 309324 326334 309376 326340
rect 309336 29646 309364 326334
rect 309324 29640 309376 29646
rect 309324 29582 309376 29588
rect 309232 28280 309284 28286
rect 309232 28222 309284 28228
rect 307116 24200 307168 24206
rect 307116 24142 307168 24148
rect 309428 17270 309456 338014
rect 309704 336530 309732 338014
rect 309692 336524 309744 336530
rect 309692 336466 309744 336472
rect 310072 326398 310100 338014
rect 310670 337770 310698 338028
rect 310808 338014 311052 338042
rect 311176 338014 311420 338042
rect 311544 338014 311788 338042
rect 311912 338014 312156 338042
rect 312280 338014 312524 338042
rect 312648 338014 312892 338042
rect 313016 338014 313260 338042
rect 313384 338014 313628 338042
rect 313752 338014 313996 338042
rect 314120 338014 314364 338042
rect 310670 337742 310744 337770
rect 310060 326392 310112 326398
rect 310060 326334 310112 326340
rect 310612 326392 310664 326398
rect 310612 326334 310664 326340
rect 310624 31074 310652 326334
rect 310716 49026 310744 337742
rect 310808 336122 310836 338014
rect 310796 336116 310848 336122
rect 310796 336058 310848 336064
rect 311176 326398 311204 338014
rect 311164 326392 311216 326398
rect 311164 326334 311216 326340
rect 311544 316034 311572 338014
rect 311912 336190 311940 338014
rect 312280 336682 312308 338014
rect 312004 336654 312308 336682
rect 311900 336184 311952 336190
rect 311900 336126 311952 336132
rect 310808 316006 311572 316034
rect 310704 49020 310756 49026
rect 310704 48962 310756 48968
rect 310704 39364 310756 39370
rect 310704 39306 310756 39312
rect 310612 31068 310664 31074
rect 310612 31010 310664 31016
rect 309416 17264 309468 17270
rect 309416 17206 309468 17212
rect 310716 16574 310744 39306
rect 310808 22846 310836 316006
rect 312004 32434 312032 336654
rect 312648 335354 312676 338014
rect 312096 335326 312676 335354
rect 312096 50386 312124 335326
rect 313016 316034 313044 338014
rect 313384 336734 313412 338014
rect 313372 336728 313424 336734
rect 313372 336670 313424 336676
rect 313752 335354 313780 338014
rect 312188 316006 313044 316034
rect 313384 335326 313780 335354
rect 313924 335368 313976 335374
rect 312084 50380 312136 50386
rect 312084 50322 312136 50328
rect 311992 32428 312044 32434
rect 311992 32370 312044 32376
rect 310796 22840 310848 22846
rect 310796 22782 310848 22788
rect 310716 16546 311480 16574
rect 307024 11824 307076 11830
rect 307024 11766 307076 11772
rect 307944 11756 307996 11762
rect 307944 11698 307996 11704
rect 306564 6316 306616 6322
rect 306564 6258 306616 6264
rect 304264 6248 304316 6254
rect 304264 6190 304316 6196
rect 306748 6180 306800 6186
rect 306748 6122 306800 6128
rect 305552 4140 305604 4146
rect 305552 4082 305604 4088
rect 305564 480 305592 4082
rect 306760 480 306788 6122
rect 307956 480 307984 11698
rect 310244 7608 310296 7614
rect 310244 7550 310296 7556
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 7550
rect 311452 480 311480 16546
rect 312188 9110 312216 316006
rect 313384 51746 313412 335326
rect 313924 335310 313976 335316
rect 313464 330540 313516 330546
rect 313464 330482 313516 330488
rect 313372 51740 313424 51746
rect 313372 51682 313424 51688
rect 313476 21486 313504 330482
rect 313464 21480 313516 21486
rect 313464 21422 313516 21428
rect 313936 14482 313964 335310
rect 314120 330546 314148 338014
rect 314718 337770 314746 338028
rect 314856 338014 315100 338042
rect 315224 338014 315468 338042
rect 315592 338014 315836 338042
rect 314718 337742 314792 337770
rect 314108 330540 314160 330546
rect 314108 330482 314160 330488
rect 314764 33794 314792 337742
rect 314856 336666 314884 338014
rect 314844 336660 314896 336666
rect 314844 336602 314896 336608
rect 315224 336054 315252 338014
rect 315304 336320 315356 336326
rect 315304 336262 315356 336268
rect 315212 336048 315264 336054
rect 315212 335990 315264 335996
rect 314844 328840 314896 328846
rect 314844 328782 314896 328788
rect 314752 33788 314804 33794
rect 314752 33730 314804 33736
rect 313924 14476 313976 14482
rect 313924 14418 313976 14424
rect 313832 14000 313884 14006
rect 313832 13942 313884 13948
rect 312176 9104 312228 9110
rect 312176 9046 312228 9052
rect 312636 3324 312688 3330
rect 312636 3266 312688 3272
rect 312648 480 312676 3266
rect 313844 480 313872 13942
rect 314856 8974 314884 328782
rect 315316 18698 315344 336262
rect 315592 328846 315620 338014
rect 316190 337770 316218 338028
rect 316328 338014 316572 338042
rect 316696 338014 316940 338042
rect 317064 338014 317308 338042
rect 317432 338014 317676 338042
rect 317800 338014 318044 338042
rect 318168 338014 318412 338042
rect 318536 338014 318780 338042
rect 318904 338014 319148 338042
rect 319272 338014 319424 338042
rect 319548 338014 319792 338042
rect 319916 338014 320160 338042
rect 320284 338014 320528 338042
rect 320652 338014 320896 338042
rect 321020 338014 321264 338042
rect 316190 337742 316264 337770
rect 316132 336728 316184 336734
rect 316132 336670 316184 336676
rect 315580 328840 315632 328846
rect 315580 328782 315632 328788
rect 316144 22778 316172 336670
rect 316236 26994 316264 337742
rect 316328 336734 316356 338014
rect 316316 336728 316368 336734
rect 316316 336670 316368 336676
rect 316696 336258 316724 338014
rect 316684 336252 316736 336258
rect 316684 336194 316736 336200
rect 317064 316034 317092 338014
rect 317432 335374 317460 338014
rect 317420 335368 317472 335374
rect 317800 335354 317828 338014
rect 318064 336116 318116 336122
rect 318064 336058 318116 336064
rect 317420 335310 317472 335316
rect 317616 335326 317828 335354
rect 317512 330472 317564 330478
rect 317512 330414 317564 330420
rect 316328 316006 317092 316034
rect 316224 26988 316276 26994
rect 316224 26930 316276 26936
rect 316132 22772 316184 22778
rect 316132 22714 316184 22720
rect 315304 18692 315356 18698
rect 315304 18634 315356 18640
rect 314844 8968 314896 8974
rect 314844 8910 314896 8916
rect 316328 3534 316356 316006
rect 317524 13122 317552 330414
rect 317616 35222 317644 335326
rect 317696 330540 317748 330546
rect 317696 330482 317748 330488
rect 317604 35216 317656 35222
rect 317604 35158 317656 35164
rect 317512 13116 317564 13122
rect 317512 13058 317564 13064
rect 317328 8968 317380 8974
rect 317328 8910 317380 8916
rect 316316 3528 316368 3534
rect 316316 3470 316368 3476
rect 316224 3460 316276 3466
rect 316224 3402 316276 3408
rect 315028 3256 315080 3262
rect 315028 3198 315080 3204
rect 315040 480 315068 3198
rect 316236 480 316264 3402
rect 317340 480 317368 8910
rect 317708 3194 317736 330482
rect 318076 14006 318104 336058
rect 318168 330546 318196 338014
rect 318156 330540 318208 330546
rect 318156 330482 318208 330488
rect 318536 330478 318564 338014
rect 318800 330540 318852 330546
rect 318800 330482 318852 330488
rect 318524 330472 318576 330478
rect 318524 330414 318576 330420
rect 318064 14000 318116 14006
rect 318064 13942 318116 13948
rect 318812 3602 318840 330482
rect 318904 7750 318932 338014
rect 319272 330546 319300 338014
rect 319548 336682 319576 338014
rect 319364 336654 319576 336682
rect 319260 330540 319312 330546
rect 319260 330482 319312 330488
rect 318984 330472 319036 330478
rect 318984 330414 319036 330420
rect 318996 250646 319024 330414
rect 319364 316034 319392 336654
rect 319444 335844 319496 335850
rect 319444 335786 319496 335792
rect 319088 316006 319392 316034
rect 319088 274106 319116 316006
rect 319076 274100 319128 274106
rect 319076 274042 319128 274048
rect 318984 250640 319036 250646
rect 318984 250582 319036 250588
rect 319456 15910 319484 335786
rect 319916 330478 319944 338014
rect 320180 336048 320232 336054
rect 320180 335990 320232 335996
rect 319904 330472 319956 330478
rect 319904 330414 319956 330420
rect 319444 15904 319496 15910
rect 319444 15846 319496 15852
rect 318892 7744 318944 7750
rect 318892 7686 318944 7692
rect 318800 3596 318852 3602
rect 318800 3538 318852 3544
rect 319720 3596 319772 3602
rect 319720 3538 319772 3544
rect 318524 3528 318576 3534
rect 318524 3470 318576 3476
rect 317696 3188 317748 3194
rect 317696 3130 317748 3136
rect 318536 480 318564 3470
rect 319732 480 319760 3538
rect 320192 490 320220 335990
rect 320284 3369 320312 338014
rect 320652 316034 320680 338014
rect 321020 335850 321048 338014
rect 321618 337770 321646 338028
rect 321756 338014 322000 338042
rect 322124 338014 322368 338042
rect 322492 338014 322736 338042
rect 321618 337742 321692 337770
rect 321008 335844 321060 335850
rect 321008 335786 321060 335792
rect 320824 335776 320876 335782
rect 320824 335718 320876 335724
rect 320376 316006 320680 316034
rect 320376 4894 320404 316006
rect 320836 279682 320864 335718
rect 321560 326392 321612 326398
rect 321560 326334 321612 326340
rect 320824 279676 320876 279682
rect 320824 279618 320876 279624
rect 320364 4888 320416 4894
rect 320364 4830 320416 4836
rect 321572 3738 321600 326334
rect 321560 3732 321612 3738
rect 321560 3674 321612 3680
rect 321664 3670 321692 337742
rect 321756 24138 321784 338014
rect 322124 316034 322152 338014
rect 322492 326398 322520 338014
rect 323090 337770 323118 338028
rect 323228 338014 323472 338042
rect 323596 338014 323840 338042
rect 323964 338014 324208 338042
rect 324332 338014 324576 338042
rect 324700 338014 324944 338042
rect 325068 338014 325312 338042
rect 325436 338014 325680 338042
rect 325896 338014 326048 338042
rect 326172 338014 326416 338042
rect 326540 338014 326784 338042
rect 323090 337742 323164 337770
rect 323032 326460 323084 326466
rect 323032 326402 323084 326408
rect 322480 326392 322532 326398
rect 322480 326334 322532 326340
rect 322940 326392 322992 326398
rect 322940 326334 322992 326340
rect 321848 316006 322152 316034
rect 321848 36582 321876 316006
rect 321836 36576 321888 36582
rect 321836 36518 321888 36524
rect 321744 24132 321796 24138
rect 321744 24074 321796 24080
rect 322952 3806 322980 326334
rect 323044 10402 323072 326402
rect 323136 25566 323164 337742
rect 323228 284986 323256 338014
rect 323596 326398 323624 338014
rect 323964 326466 323992 338014
rect 324332 336326 324360 338014
rect 324700 336682 324728 338014
rect 324424 336654 324728 336682
rect 324320 336320 324372 336326
rect 324320 336262 324372 336268
rect 324320 336184 324372 336190
rect 324320 336126 324372 336132
rect 323952 326460 324004 326466
rect 323952 326402 324004 326408
rect 323584 326392 323636 326398
rect 323584 326334 323636 326340
rect 323216 284980 323268 284986
rect 323216 284922 323268 284928
rect 323124 25560 323176 25566
rect 323124 25502 323176 25508
rect 323032 10396 323084 10402
rect 323032 10338 323084 10344
rect 322940 3800 322992 3806
rect 322940 3742 322992 3748
rect 323308 3732 323360 3738
rect 323308 3674 323360 3680
rect 321652 3664 321704 3670
rect 321652 3606 321704 3612
rect 322112 3664 322164 3670
rect 322112 3606 322164 3612
rect 320270 3360 320326 3369
rect 320270 3295 320326 3304
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320192 462 320496 490
rect 322124 480 322152 3606
rect 323320 480 323348 3674
rect 324332 3482 324360 336126
rect 324424 3874 324452 336654
rect 325068 335354 325096 338014
rect 324516 335326 325096 335354
rect 324516 4826 324544 335326
rect 325436 316034 325464 338014
rect 325896 328454 325924 338014
rect 326172 335354 326200 338014
rect 326540 335782 326568 338014
rect 327138 337770 327166 338028
rect 327276 338014 327520 338042
rect 327644 338014 327888 338042
rect 328012 338014 328256 338042
rect 328564 338014 328624 338042
rect 328748 338014 328992 338042
rect 329116 338014 329360 338042
rect 329484 338014 329728 338042
rect 330036 338014 330096 338042
rect 330220 338014 330464 338042
rect 330588 338014 330832 338042
rect 330956 338014 331108 338042
rect 331324 338014 331476 338042
rect 331600 338014 331844 338042
rect 331968 338014 332212 338042
rect 332336 338014 332580 338042
rect 332796 338014 332948 338042
rect 333072 338014 333316 338042
rect 333440 338014 333684 338042
rect 333992 338014 334052 338042
rect 334176 338014 334420 338042
rect 334544 338014 334788 338042
rect 334912 338014 335156 338042
rect 335464 338014 335524 338042
rect 335648 338014 335892 338042
rect 336016 338014 336260 338042
rect 336384 338014 336628 338042
rect 336844 338014 336996 338042
rect 337120 338014 337364 338042
rect 337488 338014 337732 338042
rect 337856 338014 338100 338042
rect 338224 338014 338468 338042
rect 338592 338014 338836 338042
rect 338960 338014 339204 338042
rect 327138 337742 327212 337770
rect 326528 335776 326580 335782
rect 326528 335718 326580 335724
rect 325804 328426 325924 328454
rect 325988 335326 326200 335354
rect 325804 323626 325832 328426
rect 325804 323598 325924 323626
rect 325792 319524 325844 319530
rect 325792 319466 325844 319472
rect 324608 316006 325464 316034
rect 324608 261594 324636 316006
rect 324596 261588 324648 261594
rect 324596 261530 324648 261536
rect 325804 4962 325832 319466
rect 325792 4956 325844 4962
rect 325792 4898 325844 4904
rect 324504 4820 324556 4826
rect 324504 4762 324556 4768
rect 325896 3942 325924 323598
rect 325988 319530 326016 335326
rect 327080 326392 327132 326398
rect 327080 326334 327132 326340
rect 325976 319524 326028 319530
rect 325976 319466 326028 319472
rect 327092 4078 327120 326334
rect 327080 4072 327132 4078
rect 327080 4014 327132 4020
rect 327184 4010 327212 337742
rect 327276 5030 327304 338014
rect 327644 316034 327672 338014
rect 328012 326398 328040 338014
rect 328460 326460 328512 326466
rect 328460 326402 328512 326408
rect 328000 326392 328052 326398
rect 328000 326334 328052 326340
rect 327368 316006 327672 316034
rect 327368 254794 327396 316006
rect 327356 254788 327408 254794
rect 327356 254730 327408 254736
rect 327264 5024 327316 5030
rect 327264 4966 327316 4972
rect 328472 4146 328500 326402
rect 328564 5098 328592 338014
rect 328644 326392 328696 326398
rect 328644 326334 328696 326340
rect 328656 6186 328684 326334
rect 328748 253434 328776 338014
rect 329116 326466 329144 338014
rect 329104 326460 329156 326466
rect 329104 326402 329156 326408
rect 329484 326398 329512 338014
rect 329932 326460 329984 326466
rect 329932 326402 329984 326408
rect 329472 326392 329524 326398
rect 329472 326334 329524 326340
rect 329840 326392 329892 326398
rect 329840 326334 329892 326340
rect 328736 253428 328788 253434
rect 328736 253370 328788 253376
rect 328644 6180 328696 6186
rect 328644 6122 328696 6128
rect 328552 5092 328604 5098
rect 328552 5034 328604 5040
rect 328460 4140 328512 4146
rect 328460 4082 328512 4088
rect 327172 4004 327224 4010
rect 327172 3946 327224 3952
rect 325884 3936 325936 3942
rect 325884 3878 325936 3884
rect 326804 3936 326856 3942
rect 326804 3878 326856 3884
rect 328000 3936 328052 3942
rect 328000 3878 328052 3884
rect 324412 3868 324464 3874
rect 324412 3810 324464 3816
rect 325608 3800 325660 3806
rect 325608 3742 325660 3748
rect 324332 3454 324452 3482
rect 324424 480 324452 3454
rect 325620 480 325648 3742
rect 326816 480 326844 3878
rect 328012 480 328040 3878
rect 329196 3868 329248 3874
rect 329196 3810 329248 3816
rect 329208 480 329236 3810
rect 329852 3398 329880 326334
rect 329944 7614 329972 326402
rect 330036 11762 330064 338014
rect 330220 326398 330248 338014
rect 330588 326466 330616 338014
rect 330576 326460 330628 326466
rect 330576 326402 330628 326408
rect 330208 326392 330260 326398
rect 330208 326334 330260 326340
rect 330956 316034 330984 338014
rect 331220 336932 331272 336938
rect 331220 336874 331272 336880
rect 331232 336122 331260 336874
rect 331220 336116 331272 336122
rect 331220 336058 331272 336064
rect 330128 316006 330984 316034
rect 330128 39370 330156 316006
rect 330116 39364 330168 39370
rect 330116 39306 330168 39312
rect 330024 11756 330076 11762
rect 330024 11698 330076 11704
rect 329932 7608 329984 7614
rect 329932 7550 329984 7556
rect 329840 3392 329892 3398
rect 329840 3334 329892 3340
rect 331324 3330 331352 338014
rect 331600 336938 331628 338014
rect 331588 336932 331640 336938
rect 331588 336874 331640 336880
rect 331968 336818 331996 338014
rect 331416 336790 331996 336818
rect 331312 3324 331364 3330
rect 331312 3266 331364 3272
rect 331416 3262 331444 336790
rect 332336 336682 332364 338014
rect 331508 336654 332364 336682
rect 331508 3466 331536 336654
rect 331588 335368 331640 335374
rect 331588 335310 331640 335316
rect 331496 3460 331548 3466
rect 331496 3402 331548 3408
rect 331404 3256 331456 3262
rect 331404 3198 331456 3204
rect 330392 3188 330444 3194
rect 330392 3130 330444 3136
rect 330404 480 330432 3130
rect 331600 480 331628 335310
rect 332600 330540 332652 330546
rect 332600 330482 332652 330488
rect 332612 4434 332640 330482
rect 332692 330472 332744 330478
rect 332692 330414 332744 330420
rect 332520 4406 332640 4434
rect 332520 3534 332548 4406
rect 332704 4298 332732 330414
rect 332796 8974 332824 338014
rect 333072 330546 333100 338014
rect 333060 330540 333112 330546
rect 333060 330482 333112 330488
rect 333440 330478 333468 338014
rect 333992 336054 334020 338014
rect 333980 336048 334032 336054
rect 333980 335990 334032 335996
rect 334176 335354 334204 338014
rect 334544 336682 334572 338014
rect 334084 335326 334204 335354
rect 334268 336654 334572 336682
rect 333428 330472 333480 330478
rect 333428 330414 333480 330420
rect 332784 8968 332836 8974
rect 332784 8910 332836 8916
rect 332612 4270 332732 4298
rect 332612 3602 332640 4270
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 332600 3596 332652 3602
rect 332600 3538 332652 3544
rect 332508 3528 332560 3534
rect 332508 3470 332560 3476
rect 332704 480 332732 4082
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 333900 480 333928 3946
rect 334084 3670 334112 335326
rect 334268 316034 334296 336654
rect 334348 336320 334400 336326
rect 334348 336262 334400 336268
rect 334176 316006 334296 316034
rect 334176 3738 334204 316006
rect 334360 16574 334388 336262
rect 334912 336190 334940 338014
rect 334900 336184 334952 336190
rect 334900 336126 334952 336132
rect 335360 330540 335412 330546
rect 335360 330482 335412 330488
rect 334360 16546 334664 16574
rect 334164 3732 334216 3738
rect 334164 3674 334216 3680
rect 334072 3664 334124 3670
rect 334072 3606 334124 3612
rect 320468 354 320496 462
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335372 3942 335400 330482
rect 335360 3936 335412 3942
rect 335360 3878 335412 3884
rect 335464 3806 335492 338014
rect 335648 335354 335676 338014
rect 335556 335326 335676 335354
rect 335556 4078 335584 335326
rect 336016 330546 336044 338014
rect 336004 330540 336056 330546
rect 336004 330482 336056 330488
rect 336384 316034 336412 338014
rect 335648 316006 336412 316034
rect 335544 4072 335596 4078
rect 335544 4014 335596 4020
rect 335648 3874 335676 316006
rect 335636 3868 335688 3874
rect 335636 3810 335688 3816
rect 335452 3800 335504 3806
rect 335452 3742 335504 3748
rect 336844 3262 336872 338014
rect 337120 335374 337148 338014
rect 337108 335368 337160 335374
rect 337488 335354 337516 338014
rect 337108 335310 337160 335316
rect 337212 335326 337516 335354
rect 337212 330528 337240 335326
rect 336936 330500 337240 330528
rect 336936 4146 336964 330500
rect 337856 316034 337884 338014
rect 338224 336326 338252 338014
rect 338212 336320 338264 336326
rect 338212 336262 338264 336268
rect 338592 335354 338620 338014
rect 338316 335326 338620 335354
rect 338316 316034 338344 335326
rect 338960 316034 338988 338014
rect 339558 337770 339586 338028
rect 339696 338014 339940 338042
rect 340064 338014 340308 338042
rect 340676 338014 340828 338042
rect 339558 337742 339632 337770
rect 339500 336252 339552 336258
rect 339500 336194 339552 336200
rect 337120 316006 337884 316034
rect 338224 316006 338344 316034
rect 338408 316006 338988 316034
rect 336924 4140 336976 4146
rect 336924 4082 336976 4088
rect 337120 4010 337148 316006
rect 337108 4004 337160 4010
rect 337108 3946 337160 3952
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 336832 3256 336884 3262
rect 336832 3198 336884 3204
rect 336280 3188 336332 3194
rect 336280 3130 336332 3136
rect 336292 480 336320 3130
rect 337488 480 337516 3470
rect 338224 3194 338252 316006
rect 338408 3534 338436 316006
rect 338396 3528 338448 3534
rect 338396 3470 338448 3476
rect 338672 3528 338724 3534
rect 338672 3470 338724 3476
rect 338212 3188 338264 3194
rect 338212 3130 338264 3136
rect 338684 480 338712 3470
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 336194
rect 339604 3534 339632 337742
rect 339696 336258 339724 338014
rect 339684 336252 339736 336258
rect 339684 336194 339736 336200
rect 340064 316034 340092 338014
rect 340800 336598 340828 338014
rect 340984 338014 341044 338042
rect 341168 338014 341412 338042
rect 341536 338014 341780 338042
rect 341904 338014 342148 338042
rect 340788 336592 340840 336598
rect 340788 336534 340840 336540
rect 340984 335714 341012 338014
rect 340972 335708 341024 335714
rect 340972 335650 341024 335656
rect 341168 335354 341196 338014
rect 341536 336682 341564 338014
rect 341076 335326 341196 335354
rect 341260 336654 341564 336682
rect 340972 326392 341024 326398
rect 340972 326334 341024 326340
rect 339696 316006 340092 316034
rect 339696 3534 339724 316006
rect 340984 4078 341012 326334
rect 340972 4072 341024 4078
rect 340972 4014 341024 4020
rect 339592 3528 339644 3534
rect 339592 3470 339644 3476
rect 339684 3528 339736 3534
rect 339684 3470 339736 3476
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 340984 480 341012 3470
rect 341076 3398 341104 335326
rect 341260 316034 341288 336654
rect 341340 336592 341392 336598
rect 341340 336534 341392 336540
rect 341168 316006 341288 316034
rect 341168 4146 341196 316006
rect 341352 16574 341380 336534
rect 341904 326398 341932 338014
rect 342502 337770 342530 338028
rect 342640 338014 342884 338042
rect 343008 338014 343160 338042
rect 343284 338014 343528 338042
rect 343836 338014 343896 338042
rect 344020 338014 344264 338042
rect 344388 338014 344632 338042
rect 344940 338014 345000 338042
rect 345124 338014 345368 338042
rect 345676 338014 345736 338042
rect 345860 338014 346104 338042
rect 346472 338014 346624 338042
rect 342502 337742 342576 337770
rect 342444 336728 342496 336734
rect 342444 336670 342496 336676
rect 342260 335708 342312 335714
rect 342260 335650 342312 335656
rect 341892 326392 341944 326398
rect 341892 326334 341944 326340
rect 341352 16546 342208 16574
rect 341156 4140 341208 4146
rect 341156 4082 341208 4088
rect 341064 3392 341116 3398
rect 341064 3334 341116 3340
rect 342180 480 342208 16546
rect 342272 2530 342300 335650
rect 342352 326392 342404 326398
rect 342352 326334 342404 326340
rect 342364 3602 342392 326334
rect 342456 3738 342484 336670
rect 342548 3942 342576 337742
rect 342640 336734 342668 338014
rect 342628 336728 342680 336734
rect 342628 336670 342680 336676
rect 343008 316034 343036 338014
rect 343284 326398 343312 338014
rect 343836 336190 343864 338014
rect 343824 336184 343876 336190
rect 343824 336126 343876 336132
rect 343272 326392 343324 326398
rect 343272 326334 343324 326340
rect 343640 323332 343692 323338
rect 343640 323274 343692 323280
rect 342640 316006 343036 316034
rect 342536 3936 342588 3942
rect 342536 3878 342588 3884
rect 342640 3874 342668 316006
rect 342628 3868 342680 3874
rect 342628 3810 342680 3816
rect 342444 3732 342496 3738
rect 342444 3674 342496 3680
rect 342352 3596 342404 3602
rect 342352 3538 342404 3544
rect 343652 3466 343680 323274
rect 344020 316034 344048 338014
rect 344388 323338 344416 338014
rect 344940 336054 344968 338014
rect 344928 336048 344980 336054
rect 344928 335990 344980 335996
rect 344376 323332 344428 323338
rect 344376 323274 344428 323280
rect 345020 322244 345072 322250
rect 345020 322186 345072 322192
rect 343744 316006 344048 316034
rect 343744 3534 343772 316006
rect 345032 6254 345060 322186
rect 345124 10402 345152 338014
rect 345676 336326 345704 338014
rect 345664 336320 345716 336326
rect 345664 336262 345716 336268
rect 345664 336184 345716 336190
rect 345664 336126 345716 336132
rect 345112 10396 345164 10402
rect 345112 10338 345164 10344
rect 345020 6248 345072 6254
rect 345020 6190 345072 6196
rect 345676 4214 345704 336126
rect 345860 322250 345888 338014
rect 346400 336728 346452 336734
rect 346400 336670 346452 336676
rect 345848 322244 345900 322250
rect 345848 322186 345900 322192
rect 345664 4208 345716 4214
rect 345664 4150 345716 4156
rect 345756 4140 345808 4146
rect 345756 4082 345808 4088
rect 343732 3528 343784 3534
rect 343732 3470 343784 3476
rect 343640 3460 343692 3466
rect 343640 3402 343692 3408
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 342272 2502 342944 2530
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 2502
rect 344572 480 344600 3334
rect 345768 480 345796 4082
rect 346412 3670 346440 336670
rect 346492 326392 346544 326398
rect 346492 326334 346544 326340
rect 346504 6186 346532 326334
rect 346596 17270 346624 338014
rect 346688 338014 346840 338042
rect 347208 338014 347360 338042
rect 346688 336734 346716 338014
rect 346676 336728 346728 336734
rect 346676 336670 346728 336676
rect 347332 336258 347360 338014
rect 347424 338014 347576 338042
rect 347320 336252 347372 336258
rect 347320 336194 347372 336200
rect 347424 326398 347452 338014
rect 347930 337770 347958 338028
rect 348068 338014 348312 338042
rect 348620 338014 348680 338042
rect 348804 338014 349048 338042
rect 349172 338014 349416 338042
rect 349540 338014 349784 338042
rect 350092 338014 350152 338042
rect 350276 338014 350520 338042
rect 350828 338014 350888 338042
rect 351012 338014 351256 338042
rect 351380 338014 351624 338042
rect 351932 338014 351992 338042
rect 352116 338014 352360 338042
rect 352484 338014 352728 338042
rect 352852 338014 353096 338042
rect 353312 338014 353464 338042
rect 353772 338014 353832 338042
rect 353956 338014 354200 338042
rect 354324 338014 354568 338042
rect 347930 337742 348004 337770
rect 347976 328454 348004 337742
rect 347884 328426 348004 328454
rect 347412 326392 347464 326398
rect 347412 326334 347464 326340
rect 347780 323876 347832 323882
rect 347780 323818 347832 323824
rect 346584 17264 346636 17270
rect 346584 17206 346636 17212
rect 347792 7614 347820 323818
rect 347884 321858 347912 328426
rect 347884 321830 348004 321858
rect 347872 321564 347924 321570
rect 347872 321506 347924 321512
rect 347884 7682 347912 321506
rect 347976 26926 348004 321830
rect 348068 321570 348096 338014
rect 348620 336190 348648 338014
rect 348608 336184 348660 336190
rect 348608 336126 348660 336132
rect 348804 323882 348832 338014
rect 348792 323876 348844 323882
rect 348792 323818 348844 323824
rect 348056 321564 348108 321570
rect 348056 321506 348108 321512
rect 347964 26920 348016 26926
rect 347964 26862 348016 26868
rect 349172 9042 349200 338014
rect 349540 335354 349568 338014
rect 350092 336530 350120 338014
rect 350080 336524 350132 336530
rect 350080 336466 350132 336472
rect 349264 335326 349568 335354
rect 349264 10334 349292 335326
rect 350276 316034 350304 338014
rect 350828 336122 350856 338014
rect 350816 336116 350868 336122
rect 350816 336058 350868 336064
rect 350540 326392 350592 326398
rect 350540 326334 350592 326340
rect 349356 316006 350304 316034
rect 349356 11830 349384 316006
rect 350552 13190 350580 326334
rect 351012 316034 351040 338014
rect 351184 336048 351236 336054
rect 351184 335990 351236 335996
rect 350644 316006 351040 316034
rect 350644 28286 350672 316006
rect 350632 28280 350684 28286
rect 350632 28222 350684 28228
rect 350540 13184 350592 13190
rect 350540 13126 350592 13132
rect 349344 11824 349396 11830
rect 349344 11766 349396 11772
rect 349252 10328 349304 10334
rect 349252 10270 349304 10276
rect 349160 9036 349212 9042
rect 349160 8978 349212 8984
rect 347872 7676 347924 7682
rect 347872 7618 347924 7624
rect 347780 7608 347832 7614
rect 347780 7550 347832 7556
rect 346492 6180 346544 6186
rect 346492 6122 346544 6128
rect 351196 4962 351224 335990
rect 351380 326398 351408 338014
rect 351932 336054 351960 338014
rect 351920 336048 351972 336054
rect 351920 335990 351972 335996
rect 352116 335866 352144 338014
rect 351932 335838 352144 335866
rect 351368 326392 351420 326398
rect 351368 326334 351420 326340
rect 351932 8974 351960 335838
rect 352484 335354 352512 338014
rect 352024 335326 352512 335354
rect 352024 14482 352052 335326
rect 352852 316034 352880 338014
rect 352116 316006 352880 316034
rect 352116 21418 352144 316006
rect 352104 21412 352156 21418
rect 352104 21354 352156 21360
rect 352012 14476 352064 14482
rect 352012 14418 352064 14424
rect 351920 8968 351972 8974
rect 351920 8910 351972 8916
rect 351184 4956 351236 4962
rect 351184 4898 351236 4904
rect 353312 4894 353340 338014
rect 353772 336462 353800 338014
rect 353760 336456 353812 336462
rect 353760 336398 353812 336404
rect 353956 335354 353984 338014
rect 353404 335326 353984 335354
rect 353404 24274 353432 335326
rect 354324 316034 354352 338014
rect 354922 337770 354950 338028
rect 355060 338014 355212 338042
rect 355336 338014 355580 338042
rect 355704 338014 355948 338042
rect 356256 338014 356316 338042
rect 356440 338014 356684 338042
rect 356808 338014 357052 338042
rect 357176 338014 357420 338042
rect 357636 338014 357788 338042
rect 354922 337742 354996 337770
rect 354968 326534 354996 337742
rect 354956 326528 355008 326534
rect 354956 326470 355008 326476
rect 354680 326460 354732 326466
rect 354680 326402 354732 326408
rect 353496 316006 354352 316034
rect 353496 243574 353524 316006
rect 353484 243568 353536 243574
rect 353484 243510 353536 243516
rect 353392 24268 353444 24274
rect 353392 24210 353444 24216
rect 353300 4888 353352 4894
rect 353300 4830 353352 4836
rect 354692 4826 354720 326402
rect 354772 326392 354824 326398
rect 354772 326334 354824 326340
rect 354784 29646 354812 326334
rect 355060 323626 355088 338014
rect 355140 326528 355192 326534
rect 355140 326470 355192 326476
rect 354876 323598 355088 323626
rect 354876 261526 354904 323598
rect 355152 318794 355180 326470
rect 355336 326398 355364 338014
rect 355704 326466 355732 338014
rect 356256 326466 356284 338014
rect 356440 335354 356468 338014
rect 356348 335326 356468 335354
rect 355692 326460 355744 326466
rect 355692 326402 355744 326408
rect 356244 326460 356296 326466
rect 356244 326402 356296 326408
rect 355324 326392 355376 326398
rect 355324 326334 355376 326340
rect 356060 326392 356112 326398
rect 356060 326334 356112 326340
rect 354968 318766 355180 318794
rect 354968 286414 354996 318766
rect 354956 286408 355008 286414
rect 354956 286350 355008 286356
rect 354864 261520 354916 261526
rect 354864 261462 354916 261468
rect 354772 29640 354824 29646
rect 354772 29582 354824 29588
rect 356072 22778 356100 326334
rect 356348 323626 356376 335326
rect 356428 326460 356480 326466
rect 356428 326402 356480 326408
rect 356164 323598 356376 323626
rect 356164 31074 356192 323598
rect 356440 318794 356468 326402
rect 356256 318766 356468 318794
rect 356256 260166 356284 318766
rect 356808 316034 356836 338014
rect 357176 326398 357204 338014
rect 357440 336320 357492 336326
rect 357440 336262 357492 336268
rect 357164 326392 357216 326398
rect 357164 326334 357216 326340
rect 356348 316006 356836 316034
rect 356348 285054 356376 316006
rect 356336 285048 356388 285054
rect 356336 284990 356388 284996
rect 356244 260160 356296 260166
rect 356244 260102 356296 260108
rect 356152 31068 356204 31074
rect 356152 31010 356204 31016
rect 356060 22772 356112 22778
rect 356060 22714 356112 22720
rect 356336 4956 356388 4962
rect 356336 4898 356388 4904
rect 354680 4820 354732 4826
rect 354680 4762 354732 4768
rect 352840 4208 352892 4214
rect 352840 4150 352892 4156
rect 346952 4072 347004 4078
rect 346952 4014 347004 4020
rect 346400 3664 346452 3670
rect 346400 3606 346452 3612
rect 346964 480 346992 4014
rect 348056 3936 348108 3942
rect 348056 3878 348108 3884
rect 348068 480 348096 3878
rect 350448 3868 350500 3874
rect 350448 3810 350500 3816
rect 349252 3732 349304 3738
rect 349252 3674 349304 3680
rect 349264 480 349292 3674
rect 350460 480 350488 3810
rect 351644 3596 351696 3602
rect 351644 3538 351696 3544
rect 351656 480 351684 3538
rect 352852 480 352880 4150
rect 354036 3528 354088 3534
rect 354036 3470 354088 3476
rect 354048 480 354076 3470
rect 355232 3460 355284 3466
rect 355232 3402 355284 3408
rect 355244 480 355272 3402
rect 356348 480 356376 4898
rect 357452 3534 357480 336262
rect 357532 326392 357584 326398
rect 357532 326334 357584 326340
rect 357544 254590 357572 326334
rect 357636 256018 357664 338014
rect 358142 337770 358170 338028
rect 358280 338014 358524 338042
rect 358892 338014 359044 338042
rect 358142 337742 358216 337770
rect 358084 336524 358136 336530
rect 358084 336466 358136 336472
rect 357624 256012 357676 256018
rect 357624 255954 357676 255960
rect 357532 254584 357584 254590
rect 357532 254526 357584 254532
rect 358096 17338 358124 336466
rect 358188 336394 358216 337742
rect 358176 336388 358228 336394
rect 358176 336330 358228 336336
rect 358280 326398 358308 338014
rect 359016 331214 359044 338014
rect 358924 331186 359044 331214
rect 359108 338014 359260 338042
rect 359384 338014 359628 338042
rect 359752 338014 359996 338042
rect 360304 338014 360364 338042
rect 360488 338014 360732 338042
rect 360856 338014 361100 338042
rect 361224 338014 361468 338042
rect 361684 338014 361836 338042
rect 361960 338014 362204 338042
rect 362572 338014 362816 338042
rect 358268 326392 358320 326398
rect 358268 326334 358320 326340
rect 358924 323626 358952 331186
rect 358820 323604 358872 323610
rect 358924 323598 359044 323626
rect 359108 323610 359136 338014
rect 358820 323546 358872 323552
rect 358084 17332 358136 17338
rect 358084 17274 358136 17280
rect 358832 15910 358860 323546
rect 358912 323264 358964 323270
rect 358912 323206 358964 323212
rect 358924 32434 358952 323206
rect 359016 253230 359044 323598
rect 359096 323604 359148 323610
rect 359096 323546 359148 323552
rect 359384 316034 359412 338014
rect 359752 323270 359780 338014
rect 360200 330540 360252 330546
rect 360200 330482 360252 330488
rect 359740 323264 359792 323270
rect 359740 323206 359792 323212
rect 359108 316006 359412 316034
rect 359108 272542 359136 316006
rect 359096 272536 359148 272542
rect 359096 272478 359148 272484
rect 359004 253224 359056 253230
rect 359004 253166 359056 253172
rect 358912 32428 358964 32434
rect 358912 32370 358964 32376
rect 358820 15904 358872 15910
rect 358820 15846 358872 15852
rect 357532 10396 357584 10402
rect 357532 10338 357584 10344
rect 357440 3528 357492 3534
rect 357440 3470 357492 3476
rect 357544 480 357572 10338
rect 359924 6248 359976 6254
rect 359924 6190 359976 6196
rect 358728 3528 358780 3534
rect 358728 3470 358780 3476
rect 358740 480 358768 3470
rect 359936 480 359964 6190
rect 360212 3602 360240 330482
rect 360304 18766 360332 338014
rect 360488 335354 360516 338014
rect 360396 335326 360516 335354
rect 360396 25566 360424 335326
rect 360856 330546 360884 338014
rect 360844 330540 360896 330546
rect 360844 330482 360896 330488
rect 361224 316034 361252 338014
rect 361580 329724 361632 329730
rect 361580 329666 361632 329672
rect 360488 316006 361252 316034
rect 360488 283694 360516 316006
rect 360476 283688 360528 283694
rect 360476 283630 360528 283636
rect 360384 25560 360436 25566
rect 360384 25502 360436 25508
rect 360292 18760 360344 18766
rect 360292 18702 360344 18708
rect 360292 17264 360344 17270
rect 360292 17206 360344 17212
rect 360304 16574 360332 17206
rect 360304 16546 361160 16574
rect 360200 3596 360252 3602
rect 360200 3538 360252 3544
rect 361132 480 361160 16546
rect 361592 3466 361620 329666
rect 361684 298790 361712 338014
rect 361960 329730 361988 338014
rect 362788 336326 362816 338014
rect 362880 338014 362940 338042
rect 363064 338014 363308 338042
rect 363432 338014 363676 338042
rect 363800 338014 364044 338042
rect 364352 338014 364412 338042
rect 364628 338014 364780 338042
rect 364904 338014 365148 338042
rect 365272 338014 365516 338042
rect 362880 336530 362908 338014
rect 362868 336524 362920 336530
rect 362868 336466 362920 336472
rect 362776 336320 362828 336326
rect 362776 336262 362828 336268
rect 362960 336252 363012 336258
rect 362960 336194 363012 336200
rect 361948 329724 362000 329730
rect 361948 329666 362000 329672
rect 361672 298784 361724 298790
rect 361672 298726 361724 298732
rect 362972 6914 363000 336194
rect 363064 13122 363092 338014
rect 363144 330540 363196 330546
rect 363144 330482 363196 330488
rect 363156 46238 363184 330482
rect 363432 316034 363460 338014
rect 363800 330546 363828 338014
rect 363788 330540 363840 330546
rect 363788 330482 363840 330488
rect 363248 316006 363460 316034
rect 363248 282266 363276 316006
rect 363236 282260 363288 282266
rect 363236 282202 363288 282208
rect 363144 46232 363196 46238
rect 363144 46174 363196 46180
rect 363052 13116 363104 13122
rect 363052 13058 363104 13064
rect 362972 6886 363552 6914
rect 362316 3664 362368 3670
rect 362316 3606 362368 3612
rect 361580 3460 361632 3466
rect 361580 3402 361632 3408
rect 362328 480 362356 3606
rect 363524 480 363552 6886
rect 364352 3262 364380 338014
rect 364432 330540 364484 330546
rect 364432 330482 364484 330488
rect 364444 3330 364472 330482
rect 364628 326398 364656 338014
rect 364616 326392 364668 326398
rect 364616 326334 364668 326340
rect 364904 316034 364932 338014
rect 365272 330546 365300 338014
rect 365870 337770 365898 338028
rect 366008 338014 366252 338042
rect 366376 338014 366620 338042
rect 366744 338014 366988 338042
rect 367264 338014 367416 338042
rect 365870 337742 365944 337770
rect 365260 330540 365312 330546
rect 365260 330482 365312 330488
rect 365812 330540 365864 330546
rect 365812 330482 365864 330488
rect 365720 327888 365772 327894
rect 365720 327830 365772 327836
rect 364536 316006 364932 316034
rect 364536 258738 364564 316006
rect 364524 258732 364576 258738
rect 364524 258674 364576 258680
rect 364616 6180 364668 6186
rect 364616 6122 364668 6128
rect 364432 3324 364484 3330
rect 364432 3266 364484 3272
rect 364340 3256 364392 3262
rect 364340 3198 364392 3204
rect 364628 480 364656 6122
rect 365732 3398 365760 327830
rect 365824 279546 365852 330482
rect 365916 280906 365944 337742
rect 366008 324970 366036 338014
rect 366272 336184 366324 336190
rect 366272 336126 366324 336132
rect 366284 325694 366312 336126
rect 366376 327894 366404 338014
rect 366744 330546 366772 338014
rect 367100 336728 367152 336734
rect 367100 336670 367152 336676
rect 366732 330540 366784 330546
rect 366732 330482 366784 330488
rect 366364 327888 366416 327894
rect 366364 327830 366416 327836
rect 366284 325666 366404 325694
rect 365996 324964 366048 324970
rect 365996 324906 366048 324912
rect 365904 280900 365956 280906
rect 365904 280842 365956 280848
rect 365812 279540 365864 279546
rect 365812 279482 365864 279488
rect 365812 26920 365864 26926
rect 365812 26862 365864 26868
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 26862
rect 366376 5574 366404 325666
rect 367008 7676 367060 7682
rect 367008 7618 367060 7624
rect 366364 5568 366416 5574
rect 366364 5510 366416 5516
rect 367020 480 367048 7618
rect 367112 4146 367140 336670
rect 367284 329112 367336 329118
rect 367284 329054 367336 329060
rect 367192 327684 367244 327690
rect 367192 327626 367244 327632
rect 367204 6526 367232 327626
rect 367296 247722 367324 329054
rect 367388 320958 367416 338014
rect 367480 338014 367632 338042
rect 367756 338014 368000 338042
rect 368124 338014 368368 338042
rect 368584 338014 368736 338042
rect 368860 338014 369104 338042
rect 369228 338014 369472 338042
rect 369596 338014 369840 338042
rect 369964 338014 370208 338042
rect 370332 338014 370576 338042
rect 370700 338014 370944 338042
rect 367480 336734 367508 338014
rect 367468 336728 367520 336734
rect 367468 336670 367520 336676
rect 367756 327690 367784 338014
rect 368124 329118 368152 338014
rect 368480 330540 368532 330546
rect 368480 330482 368532 330488
rect 368112 329112 368164 329118
rect 368112 329054 368164 329060
rect 367744 327684 367796 327690
rect 367744 327626 367796 327632
rect 367376 320952 367428 320958
rect 367376 320894 367428 320900
rect 367284 247716 367336 247722
rect 367284 247658 367336 247664
rect 367192 6520 367244 6526
rect 367192 6462 367244 6468
rect 368204 5568 368256 5574
rect 368204 5510 368256 5516
rect 367100 4140 367152 4146
rect 367100 4082 367152 4088
rect 368216 480 368244 5510
rect 368492 4010 368520 330482
rect 368584 4078 368612 338014
rect 368860 335354 368888 338014
rect 368676 335326 368888 335354
rect 368676 6458 368704 335326
rect 369228 319530 369256 338014
rect 369596 330546 369624 338014
rect 369584 330540 369636 330546
rect 369584 330482 369636 330488
rect 369860 326460 369912 326466
rect 369860 326402 369912 326408
rect 369216 319524 369268 319530
rect 369216 319466 369268 319472
rect 369400 7608 369452 7614
rect 369400 7550 369452 7556
rect 368664 6452 368716 6458
rect 368664 6394 368716 6400
rect 368572 4072 368624 4078
rect 368572 4014 368624 4020
rect 368480 4004 368532 4010
rect 368480 3946 368532 3952
rect 369412 480 369440 7550
rect 369872 3942 369900 326402
rect 369964 6390 369992 338014
rect 370332 316034 370360 338014
rect 370504 336320 370556 336326
rect 370504 336262 370556 336268
rect 370056 316006 370360 316034
rect 370056 312594 370084 316006
rect 370044 312588 370096 312594
rect 370044 312530 370096 312536
rect 370516 17270 370544 336262
rect 370700 326466 370728 338014
rect 371298 337770 371326 338028
rect 371528 338014 371680 338042
rect 371804 338014 372048 338042
rect 372172 338014 372416 338042
rect 372632 338014 372784 338042
rect 373092 338014 373152 338042
rect 373276 338014 373520 338042
rect 373644 338014 373888 338042
rect 374104 338014 374256 338042
rect 374380 338014 374624 338042
rect 374748 338014 374992 338042
rect 375300 338014 375360 338042
rect 375576 338014 375728 338042
rect 375852 338014 376096 338042
rect 376220 338014 376464 338042
rect 371298 337742 371372 337770
rect 370688 326460 370740 326466
rect 370688 326402 370740 326408
rect 371240 326324 371292 326330
rect 371240 326266 371292 326272
rect 370504 17264 370556 17270
rect 370504 17206 370556 17212
rect 370596 9036 370648 9042
rect 370596 8978 370648 8984
rect 369952 6384 370004 6390
rect 369952 6326 370004 6332
rect 369860 3936 369912 3942
rect 369860 3878 369912 3884
rect 370608 480 370636 8978
rect 371252 3874 371280 326266
rect 371344 6322 371372 337742
rect 371424 326460 371476 326466
rect 371424 326402 371476 326408
rect 371332 6316 371384 6322
rect 371332 6258 371384 6264
rect 371436 6254 371464 326402
rect 371528 318170 371556 338014
rect 371804 326330 371832 338014
rect 372172 326466 372200 338014
rect 372160 326460 372212 326466
rect 372160 326402 372212 326408
rect 371792 326324 371844 326330
rect 371792 326266 371844 326272
rect 371516 318164 371568 318170
rect 371516 318106 371568 318112
rect 372632 10878 372660 338014
rect 373092 336326 373120 338014
rect 373080 336320 373132 336326
rect 373080 336262 373132 336268
rect 373276 335354 373304 338014
rect 373356 336524 373408 336530
rect 373356 336466 373408 336472
rect 373184 335326 373304 335354
rect 372712 326460 372764 326466
rect 372712 326402 372764 326408
rect 372620 10872 372672 10878
rect 372620 10814 372672 10820
rect 372724 10810 372752 326402
rect 373184 316034 373212 335326
rect 373368 316034 373396 336466
rect 373644 326466 373672 338014
rect 374000 336116 374052 336122
rect 374000 336058 374052 336064
rect 373632 326460 373684 326466
rect 373632 326402 373684 326408
rect 372816 316006 373212 316034
rect 373276 316006 373396 316034
rect 372816 278118 372844 316006
rect 372804 278112 372856 278118
rect 372804 278054 372856 278060
rect 372804 17332 372856 17338
rect 372804 17274 372856 17280
rect 372816 16574 372844 17274
rect 372816 16546 372936 16574
rect 372712 10804 372764 10810
rect 372712 10746 372764 10752
rect 371516 10328 371568 10334
rect 371516 10270 371568 10276
rect 371424 6248 371476 6254
rect 371424 6190 371476 6196
rect 371240 3868 371292 3874
rect 371240 3810 371292 3816
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371528 354 371556 10270
rect 372908 480 372936 16546
rect 373276 11762 373304 316006
rect 373264 11756 373316 11762
rect 373264 11698 373316 11704
rect 374012 3534 374040 336058
rect 374104 6914 374132 338014
rect 374184 326460 374236 326466
rect 374184 326402 374236 326408
rect 374196 10742 374224 326402
rect 374380 316034 374408 338014
rect 374748 326466 374776 338014
rect 375300 336258 375328 338014
rect 375288 336252 375340 336258
rect 375288 336194 375340 336200
rect 375576 326534 375604 338014
rect 375852 335354 375880 338014
rect 375668 335326 375880 335354
rect 375564 326528 375616 326534
rect 375564 326470 375616 326476
rect 374736 326460 374788 326466
rect 374736 326402 374788 326408
rect 375380 326460 375432 326466
rect 375380 326402 375432 326408
rect 374288 316006 374408 316034
rect 374288 276690 374316 316006
rect 374276 276684 374328 276690
rect 374276 276626 374328 276632
rect 374276 11824 374328 11830
rect 374276 11766 374328 11772
rect 374184 10736 374236 10742
rect 374184 10678 374236 10684
rect 374104 6886 374224 6914
rect 374196 3806 374224 6886
rect 374184 3800 374236 3806
rect 374184 3742 374236 3748
rect 374000 3528 374052 3534
rect 374288 3482 374316 11766
rect 375392 3738 375420 326402
rect 375668 323626 375696 335326
rect 375748 326528 375800 326534
rect 375748 326470 375800 326476
rect 375484 323598 375696 323626
rect 375484 10674 375512 323598
rect 375760 318794 375788 326470
rect 376220 326466 376248 338014
rect 376818 337770 376846 338028
rect 376956 338014 377200 338042
rect 377324 338014 377568 338042
rect 377692 338014 377936 338042
rect 376818 337742 376892 337770
rect 376864 326466 376892 337742
rect 376208 326460 376260 326466
rect 376208 326402 376260 326408
rect 376852 326460 376904 326466
rect 376852 326402 376904 326408
rect 376956 323626 376984 338014
rect 377324 336818 377352 338014
rect 377232 336790 377352 336818
rect 377232 336190 377260 336790
rect 377692 336682 377720 338014
rect 378290 337770 378318 338028
rect 378428 338014 378672 338042
rect 378796 338014 379040 338042
rect 379164 338014 379316 338042
rect 379684 338014 379928 338042
rect 378290 337742 378364 337770
rect 377324 336654 377720 336682
rect 377220 336184 377272 336190
rect 377220 336126 377272 336132
rect 377036 326460 377088 326466
rect 377036 326402 377088 326408
rect 375576 318766 375788 318794
rect 376772 323598 376984 323626
rect 375576 275330 375604 318766
rect 375564 275324 375616 275330
rect 375564 275266 375616 275272
rect 375564 28280 375616 28286
rect 375564 28222 375616 28228
rect 375576 16574 375604 28222
rect 375576 16546 376064 16574
rect 375472 10668 375524 10674
rect 375472 10610 375524 10616
rect 375380 3732 375432 3738
rect 375380 3674 375432 3680
rect 374000 3470 374052 3476
rect 374104 3454 374316 3482
rect 375288 3528 375340 3534
rect 375288 3470 375340 3476
rect 374104 480 374132 3454
rect 375300 480 375328 3470
rect 371670 354 371782 480
rect 371528 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 376772 10606 376800 323598
rect 377048 318794 377076 326402
rect 376864 318766 377076 318794
rect 376864 273970 376892 318766
rect 377324 316034 377352 336654
rect 377404 336048 377456 336054
rect 377404 335990 377456 335996
rect 376956 316006 377352 316034
rect 376956 286346 376984 316006
rect 376944 286340 376996 286346
rect 376944 286282 376996 286288
rect 376852 273964 376904 273970
rect 376852 273906 376904 273912
rect 377312 13184 377364 13190
rect 377312 13126 377364 13132
rect 376760 10600 376812 10606
rect 376760 10542 376812 10548
rect 377324 3482 377352 13126
rect 377416 8294 377444 335990
rect 378336 326738 378364 337742
rect 378324 326732 378376 326738
rect 378324 326674 378376 326680
rect 378324 326528 378376 326534
rect 378324 326470 378376 326476
rect 378232 326324 378284 326330
rect 378232 326266 378284 326272
rect 378140 323604 378192 323610
rect 378140 323546 378192 323552
rect 377404 8288 377456 8294
rect 377404 8230 377456 8236
rect 378152 3670 378180 323546
rect 378244 10470 378272 326266
rect 378336 10538 378364 326470
rect 378428 323610 378456 338014
rect 378416 323604 378468 323610
rect 378416 323546 378468 323552
rect 378796 316034 378824 338014
rect 379164 326330 379192 338014
rect 379900 336122 379928 338014
rect 379992 338014 380052 338042
rect 380176 338014 380420 338042
rect 380544 338014 380788 338042
rect 381096 338014 381156 338042
rect 381280 338014 381524 338042
rect 381832 338014 381892 338042
rect 382016 338014 382260 338042
rect 382384 338014 382628 338042
rect 382752 338014 382996 338042
rect 383364 338014 383608 338042
rect 379888 336116 379940 336122
rect 379888 336058 379940 336064
rect 379992 335442 380020 338014
rect 379980 335436 380032 335442
rect 379980 335378 380032 335384
rect 379520 326460 379572 326466
rect 379520 326402 379572 326408
rect 379152 326324 379204 326330
rect 379152 326266 379204 326272
rect 378428 316006 378824 316034
rect 378428 284986 378456 316006
rect 378416 284980 378468 284986
rect 378416 284922 378468 284928
rect 378324 10532 378376 10538
rect 378324 10474 378376 10480
rect 378232 10464 378284 10470
rect 378232 10406 378284 10412
rect 378876 8288 378928 8294
rect 378876 8230 378928 8236
rect 378140 3664 378192 3670
rect 378140 3606 378192 3612
rect 377324 3454 377720 3482
rect 377692 480 377720 3454
rect 378888 480 378916 8230
rect 379532 3534 379560 326402
rect 380176 316034 380204 338014
rect 380544 326466 380572 338014
rect 381096 326534 381124 338014
rect 381280 335354 381308 338014
rect 381832 336054 381860 338014
rect 381820 336048 381872 336054
rect 381820 335990 381872 335996
rect 381544 335436 381596 335442
rect 381544 335378 381596 335384
rect 381188 335326 381308 335354
rect 381084 326528 381136 326534
rect 381084 326470 381136 326476
rect 380532 326460 380584 326466
rect 380532 326402 380584 326408
rect 380900 326460 380952 326466
rect 380900 326402 380952 326408
rect 379624 316006 380204 316034
rect 379624 305726 379652 316006
rect 379612 305720 379664 305726
rect 379612 305662 379664 305668
rect 379980 8968 380032 8974
rect 379980 8910 380032 8916
rect 379520 3528 379572 3534
rect 379520 3470 379572 3476
rect 379992 480 380020 8910
rect 380912 7614 380940 326402
rect 381188 323626 381216 335326
rect 381268 326528 381320 326534
rect 381268 326470 381320 326476
rect 381004 323598 381216 323626
rect 381004 10402 381032 323598
rect 381280 318794 381308 326470
rect 381096 318766 381308 318794
rect 381096 307086 381124 318766
rect 381084 307080 381136 307086
rect 381084 307022 381136 307028
rect 381556 271182 381584 335378
rect 382016 326466 382044 338014
rect 382004 326460 382056 326466
rect 382004 326402 382056 326408
rect 381544 271176 381596 271182
rect 381544 271118 381596 271124
rect 381176 14476 381228 14482
rect 381176 14418 381228 14424
rect 380992 10396 381044 10402
rect 380992 10338 381044 10344
rect 380900 7608 380952 7614
rect 380900 7550 380952 7556
rect 381188 480 381216 14418
rect 382384 10334 382412 338014
rect 382752 316034 382780 338014
rect 383014 336832 383070 336841
rect 383014 336767 383070 336776
rect 382924 336456 382976 336462
rect 382924 336398 382976 336404
rect 382568 316006 382780 316034
rect 382464 21412 382516 21418
rect 382464 21354 382516 21360
rect 382372 10328 382424 10334
rect 382372 10270 382424 10276
rect 382476 6914 382504 21354
rect 382384 6886 382504 6914
rect 382384 480 382412 6886
rect 382568 3505 382596 316006
rect 382936 4554 382964 336398
rect 383028 306338 383056 336767
rect 383580 334694 383608 338014
rect 383718 337770 383746 338028
rect 383948 338014 384100 338042
rect 383718 337742 383792 337770
rect 383568 334688 383620 334694
rect 383568 334630 383620 334636
rect 383764 326738 383792 337742
rect 383752 326732 383804 326738
rect 383752 326674 383804 326680
rect 383948 326618 383976 338014
rect 384454 337770 384482 338028
rect 384592 338014 384836 338042
rect 385144 338014 385204 338042
rect 385328 338014 385572 338042
rect 385696 338014 385940 338042
rect 386064 338014 386308 338042
rect 384454 337742 384528 337770
rect 384500 333334 384528 337742
rect 384488 333328 384540 333334
rect 384488 333270 384540 333276
rect 383672 326590 383976 326618
rect 383016 306332 383068 306338
rect 383016 306274 383068 306280
rect 383672 21418 383700 326590
rect 383844 326528 383896 326534
rect 383844 326470 383896 326476
rect 383752 326460 383804 326466
rect 383752 326402 383804 326408
rect 383764 268394 383792 326402
rect 383856 269822 383884 326470
rect 384592 326466 384620 338014
rect 384580 326460 384632 326466
rect 384580 326402 384632 326408
rect 385040 323740 385092 323746
rect 385040 323682 385092 323688
rect 383844 269816 383896 269822
rect 383844 269758 383896 269764
rect 383752 268388 383804 268394
rect 383752 268330 383804 268336
rect 385052 24138 385080 323682
rect 385144 246362 385172 338014
rect 385224 326460 385276 326466
rect 385224 326402 385276 326408
rect 385236 267034 385264 326402
rect 385328 320890 385356 338014
rect 385696 326466 385724 338014
rect 385684 326460 385736 326466
rect 385684 326402 385736 326408
rect 386064 323746 386092 338014
rect 386662 337770 386690 338028
rect 386800 338014 387044 338042
rect 387168 338014 387412 338042
rect 387536 338014 387780 338042
rect 387996 338014 388148 338042
rect 388272 338014 388516 338042
rect 388640 338014 388884 338042
rect 389192 338014 389252 338042
rect 389376 338014 389620 338042
rect 386662 337742 386736 337770
rect 386420 336728 386472 336734
rect 386420 336670 386472 336676
rect 386052 323740 386104 323746
rect 386052 323682 386104 323688
rect 385316 320884 385368 320890
rect 385316 320826 385368 320832
rect 385224 267028 385276 267034
rect 385224 266970 385276 266976
rect 386432 265674 386460 336670
rect 386604 326460 386656 326466
rect 386604 326402 386656 326408
rect 386512 323876 386564 323882
rect 386512 323818 386564 323824
rect 386420 265668 386472 265674
rect 386420 265610 386472 265616
rect 385132 246356 385184 246362
rect 385132 246298 385184 246304
rect 386524 243642 386552 323818
rect 386616 318102 386644 326402
rect 386708 319462 386736 337742
rect 386800 336734 386828 338014
rect 386788 336728 386840 336734
rect 386788 336670 386840 336676
rect 387064 336388 387116 336394
rect 387064 336330 387116 336336
rect 386696 319456 386748 319462
rect 386696 319398 386748 319404
rect 386604 318096 386656 318102
rect 386604 318038 386656 318044
rect 386512 243636 386564 243642
rect 386512 243578 386564 243584
rect 386420 243568 386472 243574
rect 386420 243510 386472 243516
rect 385132 24268 385184 24274
rect 385132 24210 385184 24216
rect 385040 24132 385092 24138
rect 385040 24074 385092 24080
rect 383660 21412 383712 21418
rect 383660 21354 383712 21360
rect 385144 16574 385172 24210
rect 386432 16574 386460 243510
rect 385144 16546 386000 16574
rect 386432 16546 386736 16574
rect 383568 4888 383620 4894
rect 383568 4830 383620 4836
rect 382924 4548 382976 4554
rect 382924 4490 382976 4496
rect 382554 3496 382610 3505
rect 382554 3431 382610 3440
rect 383580 480 383608 4830
rect 384764 4548 384816 4554
rect 384764 4490 384816 4496
rect 384776 480 384804 4490
rect 385972 480 386000 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387076 8974 387104 336330
rect 387168 323882 387196 338014
rect 387536 326466 387564 338014
rect 387524 326460 387576 326466
rect 387524 326402 387576 326408
rect 387892 326460 387944 326466
rect 387892 326402 387944 326408
rect 387800 326324 387852 326330
rect 387800 326266 387852 326272
rect 387156 323876 387208 323882
rect 387156 323818 387208 323824
rect 387812 316742 387840 326266
rect 387800 316736 387852 316742
rect 387800 316678 387852 316684
rect 387800 286408 387852 286414
rect 387800 286350 387852 286356
rect 387064 8968 387116 8974
rect 387064 8910 387116 8916
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 286350
rect 387904 242214 387932 326402
rect 387996 264246 388024 338014
rect 388272 326466 388300 338014
rect 388260 326460 388312 326466
rect 388260 326402 388312 326408
rect 388640 326330 388668 338014
rect 388628 326324 388680 326330
rect 388628 326266 388680 326272
rect 387984 264240 388036 264246
rect 387984 264182 388036 264188
rect 389192 262886 389220 338014
rect 389376 335354 389404 338014
rect 389974 337770 390002 338028
rect 390112 338014 390356 338042
rect 390664 338014 390724 338042
rect 390848 338014 391092 338042
rect 391216 338014 391368 338042
rect 391492 338014 391736 338042
rect 389974 337742 390048 337770
rect 389284 335326 389404 335354
rect 389180 262880 389232 262886
rect 389180 262822 389232 262828
rect 389180 261520 389232 261526
rect 389180 261462 389232 261468
rect 387892 242208 387944 242214
rect 387892 242150 387944 242156
rect 389192 16574 389220 261462
rect 389284 240786 389312 335326
rect 390020 330614 390048 337742
rect 390008 330608 390060 330614
rect 390008 330550 390060 330556
rect 390112 316034 390140 338014
rect 390560 330472 390612 330478
rect 390560 330414 390612 330420
rect 389376 316006 390140 316034
rect 389376 261526 389404 316006
rect 389364 261520 389416 261526
rect 389364 261462 389416 261468
rect 389272 240780 389324 240786
rect 389272 240722 389324 240728
rect 390572 26926 390600 330414
rect 390664 239426 390692 338014
rect 390744 330540 390796 330546
rect 390744 330482 390796 330488
rect 390756 283626 390784 330482
rect 390848 305658 390876 338014
rect 391216 330546 391244 338014
rect 391204 330540 391256 330546
rect 391204 330482 391256 330488
rect 391492 330478 391520 338014
rect 392090 337770 392118 338028
rect 392228 338014 392472 338042
rect 392596 338014 392840 338042
rect 392964 338014 393208 338042
rect 393516 338014 393576 338042
rect 393700 338014 393944 338042
rect 394068 338014 394312 338042
rect 394436 338014 394680 338042
rect 394804 338014 395048 338042
rect 395172 338014 395416 338042
rect 395540 338014 395784 338042
rect 396152 338014 396304 338042
rect 392090 337742 392164 337770
rect 392032 330540 392084 330546
rect 392032 330482 392084 330488
rect 391480 330472 391532 330478
rect 391480 330414 391532 330420
rect 391940 330472 391992 330478
rect 391940 330414 391992 330420
rect 391952 313954 391980 330414
rect 391940 313948 391992 313954
rect 391940 313890 391992 313896
rect 390836 305652 390888 305658
rect 390836 305594 390888 305600
rect 390744 283620 390796 283626
rect 390744 283562 390796 283568
rect 391940 260160 391992 260166
rect 391940 260102 391992 260108
rect 390652 239420 390704 239426
rect 390652 239362 390704 239368
rect 390744 29640 390796 29646
rect 390744 29582 390796 29588
rect 390560 26920 390612 26926
rect 390560 26862 390612 26868
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390756 6914 390784 29582
rect 391952 16574 391980 260102
rect 392044 238066 392072 330482
rect 392136 329118 392164 337742
rect 392124 329112 392176 329118
rect 392124 329054 392176 329060
rect 392228 316034 392256 338014
rect 392596 330546 392624 338014
rect 392584 330540 392636 330546
rect 392584 330482 392636 330488
rect 392964 330478 392992 338014
rect 393412 330540 393464 330546
rect 393412 330482 393464 330488
rect 392952 330472 393004 330478
rect 392952 330414 393004 330420
rect 393320 327684 393372 327690
rect 393320 327626 393372 327632
rect 392136 316006 392256 316034
rect 392136 260166 392164 316006
rect 392124 260160 392176 260166
rect 392124 260102 392176 260108
rect 392032 238060 392084 238066
rect 392032 238002 392084 238008
rect 393332 28286 393360 327626
rect 393424 257378 393452 330482
rect 393516 301510 393544 338014
rect 393700 327690 393728 338014
rect 394068 327758 394096 338014
rect 394436 330546 394464 338014
rect 394424 330540 394476 330546
rect 394424 330482 394476 330488
rect 394700 330540 394752 330546
rect 394700 330482 394752 330488
rect 394056 327752 394108 327758
rect 394056 327694 394108 327700
rect 393688 327684 393740 327690
rect 393688 327626 393740 327632
rect 394712 315314 394740 330482
rect 394700 315308 394752 315314
rect 394700 315250 394752 315256
rect 393504 301504 393556 301510
rect 393504 301446 393556 301452
rect 394700 285048 394752 285054
rect 394700 284990 394752 284996
rect 393412 257372 393464 257378
rect 393412 257314 393464 257320
rect 393412 31068 393464 31074
rect 393412 31010 393464 31016
rect 393320 28280 393372 28286
rect 393320 28222 393372 28228
rect 393424 16574 393452 31010
rect 394712 16574 394740 284990
rect 394804 236706 394832 338014
rect 395172 330546 395200 338014
rect 395160 330540 395212 330546
rect 395160 330482 395212 330488
rect 395540 316034 395568 338014
rect 396172 329724 396224 329730
rect 396172 329666 396224 329672
rect 396080 327820 396132 327826
rect 396080 327762 396132 327768
rect 394896 316006 395568 316034
rect 394896 282198 394924 316006
rect 394884 282192 394936 282198
rect 394884 282134 394936 282140
rect 394792 236700 394844 236706
rect 394792 236642 394844 236648
rect 396092 51746 396120 327762
rect 396184 233918 396212 329666
rect 396276 235278 396304 338014
rect 396460 338014 396520 338042
rect 396644 338014 396888 338042
rect 397012 338014 397256 338042
rect 397564 338014 397624 338042
rect 397748 338014 397992 338042
rect 398116 338014 398360 338042
rect 398484 338014 398728 338042
rect 399036 338014 399096 338042
rect 399220 338014 399464 338042
rect 399588 338014 399832 338042
rect 399956 338014 400200 338042
rect 400324 338014 400568 338042
rect 400692 338014 400936 338042
rect 401060 338014 401304 338042
rect 401672 338014 401824 338042
rect 396460 336394 396488 338014
rect 396448 336388 396500 336394
rect 396448 336330 396500 336336
rect 396644 327826 396672 338014
rect 397012 329730 397040 338014
rect 397564 331906 397592 338014
rect 397748 335354 397776 338014
rect 397656 335326 397776 335354
rect 397552 331900 397604 331906
rect 397552 331842 397604 331848
rect 397460 330540 397512 330546
rect 397656 330528 397684 335326
rect 398116 330546 398144 338014
rect 397460 330482 397512 330488
rect 397564 330500 397684 330528
rect 398104 330540 398156 330546
rect 397000 329724 397052 329730
rect 397000 329666 397052 329672
rect 396632 327820 396684 327826
rect 396632 327762 396684 327768
rect 397472 287706 397500 330482
rect 397564 300150 397592 330500
rect 398104 330482 398156 330488
rect 398484 323610 398512 338014
rect 399036 336802 399064 338014
rect 399024 336796 399076 336802
rect 399024 336738 399076 336744
rect 399220 336682 399248 338014
rect 398852 336654 399248 336682
rect 398472 323604 398524 323610
rect 398472 323546 398524 323552
rect 397552 300144 397604 300150
rect 397552 300086 397604 300092
rect 397460 287700 397512 287706
rect 397460 287642 397512 287648
rect 397460 256012 397512 256018
rect 397460 255954 397512 255960
rect 396264 235272 396316 235278
rect 396264 235214 396316 235220
rect 396172 233912 396224 233918
rect 396172 233854 396224 233860
rect 396080 51740 396132 51746
rect 396080 51682 396132 51688
rect 396080 22772 396132 22778
rect 396080 22714 396132 22720
rect 391952 16546 392624 16574
rect 393424 16546 394280 16574
rect 394712 16546 395384 16574
rect 390664 6886 390784 6914
rect 390664 480 390692 6886
rect 391848 4820 391900 4826
rect 391848 4762 391900 4768
rect 391860 480 391888 4762
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 22714
rect 397472 16574 397500 255954
rect 398852 22778 398880 336654
rect 399588 335354 399616 338014
rect 398944 335326 399616 335354
rect 398944 322250 398972 335326
rect 398932 322244 398984 322250
rect 398932 322186 398984 322192
rect 399956 316034 399984 338014
rect 400324 336682 400352 338014
rect 399036 316006 399984 316034
rect 400232 336654 400352 336682
rect 399036 254590 399064 316006
rect 398932 254584 398984 254590
rect 398932 254526 398984 254532
rect 399024 254584 399076 254590
rect 399024 254526 399076 254532
rect 398840 22772 398892 22778
rect 398840 22714 398892 22720
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398840 8968 398892 8974
rect 398840 8910 398892 8916
rect 398852 3074 398880 8910
rect 398944 3194 398972 254526
rect 400232 29646 400260 336654
rect 400692 335354 400720 338014
rect 401060 336682 401088 338014
rect 400324 335326 400720 335354
rect 400784 336654 401088 336682
rect 401600 336728 401652 336734
rect 401600 336670 401652 336676
rect 400324 311166 400352 335326
rect 400784 316034 400812 336654
rect 400864 336592 400916 336598
rect 400864 336534 400916 336540
rect 400416 316006 400812 316034
rect 400312 311160 400364 311166
rect 400312 311102 400364 311108
rect 400416 253230 400444 316006
rect 400876 256018 400904 336534
rect 400864 256012 400916 256018
rect 400864 255954 400916 255960
rect 400312 253224 400364 253230
rect 400312 253166 400364 253172
rect 400404 253224 400456 253230
rect 400404 253166 400456 253172
rect 400220 29640 400272 29646
rect 400220 29582 400272 29588
rect 400324 16574 400352 253166
rect 400324 16546 400904 16574
rect 398932 3188 398984 3194
rect 398932 3130 398984 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 401612 4826 401640 336670
rect 401692 326460 401744 326466
rect 401692 326402 401744 326408
rect 401704 229770 401732 326402
rect 401796 231130 401824 338014
rect 401888 338014 402040 338042
rect 402348 338014 402408 338042
rect 402532 338014 402776 338042
rect 403144 338014 403296 338042
rect 401888 336734 401916 338014
rect 401876 336728 401928 336734
rect 401876 336670 401928 336676
rect 402348 336462 402376 338014
rect 402336 336456 402388 336462
rect 402336 336398 402388 336404
rect 402532 326466 402560 338014
rect 402520 326460 402572 326466
rect 402520 326402 402572 326408
rect 403072 326460 403124 326466
rect 403072 326402 403124 326408
rect 402980 326324 403032 326330
rect 402980 326266 403032 326272
rect 402992 296002 403020 326266
rect 402980 295996 403032 296002
rect 402980 295938 403032 295944
rect 402980 272536 403032 272542
rect 402980 272478 403032 272484
rect 401784 231124 401836 231130
rect 401784 231066 401836 231072
rect 401692 229764 401744 229770
rect 401692 229706 401744 229712
rect 402992 16574 403020 272478
rect 403084 228410 403112 326402
rect 403164 322516 403216 322522
rect 403164 322458 403216 322464
rect 403176 251870 403204 322458
rect 403268 297430 403296 338014
rect 403360 338014 403420 338042
rect 403544 338014 403788 338042
rect 403912 338014 404156 338042
rect 404464 338014 404524 338042
rect 404648 338014 404892 338042
rect 403360 322522 403388 338014
rect 403544 326466 403572 338014
rect 403532 326460 403584 326466
rect 403532 326402 403584 326408
rect 403912 326330 403940 338014
rect 404464 326466 404492 338014
rect 404648 335354 404676 338014
rect 405246 337770 405274 338028
rect 405384 338014 405628 338042
rect 405844 338014 405996 338042
rect 406120 338014 406364 338042
rect 406488 338014 406732 338042
rect 406856 338014 407100 338042
rect 407316 338014 407468 338042
rect 407592 338014 407836 338042
rect 407960 338014 408204 338042
rect 405246 337742 405320 337770
rect 404556 335326 404676 335354
rect 404452 326460 404504 326466
rect 404452 326402 404504 326408
rect 403900 326324 403952 326330
rect 403900 326266 403952 326272
rect 404556 323626 404584 335326
rect 405292 334626 405320 337742
rect 405280 334620 405332 334626
rect 405280 334562 405332 334568
rect 404636 326460 404688 326466
rect 404636 326402 404688 326408
rect 404372 323598 404584 323626
rect 403348 322516 403400 322522
rect 403348 322458 403400 322464
rect 403256 297424 403308 297430
rect 403256 297366 403308 297372
rect 403164 251864 403216 251870
rect 403164 251806 403216 251812
rect 403072 228404 403124 228410
rect 403072 228346 403124 228352
rect 402992 16546 403664 16574
rect 402520 15904 402572 15910
rect 402520 15846 402572 15852
rect 401600 4820 401652 4826
rect 401600 4762 401652 4768
rect 402532 480 402560 15846
rect 403636 480 403664 16546
rect 404372 15910 404400 323598
rect 404648 318794 404676 326402
rect 404464 318766 404676 318794
rect 404464 250510 404492 318766
rect 405384 316034 405412 338014
rect 405740 326324 405792 326330
rect 405740 326266 405792 326272
rect 404556 316006 405412 316034
rect 404556 280838 404584 316006
rect 404544 280832 404596 280838
rect 404544 280774 404596 280780
rect 404452 250504 404504 250510
rect 404452 250446 404504 250452
rect 404452 32428 404504 32434
rect 404452 32370 404504 32376
rect 404360 15904 404412 15910
rect 404360 15846 404412 15852
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404464 354 404492 32370
rect 405752 18630 405780 326266
rect 405844 227050 405872 338014
rect 405924 326460 405976 326466
rect 405924 326402 405976 326408
rect 405936 279478 405964 326402
rect 406120 316034 406148 338014
rect 406488 326466 406516 338014
rect 406476 326460 406528 326466
rect 406476 326402 406528 326408
rect 406856 326330 406884 338014
rect 407120 326460 407172 326466
rect 407120 326402 407172 326408
rect 406844 326324 406896 326330
rect 406844 326266 406896 326272
rect 406028 316006 406148 316034
rect 406028 309806 406056 316006
rect 406016 309800 406068 309806
rect 406016 309742 406068 309748
rect 405924 279472 405976 279478
rect 405924 279414 405976 279420
rect 405832 227044 405884 227050
rect 405832 226986 405884 226992
rect 405832 18760 405884 18766
rect 405832 18702 405884 18708
rect 405740 18624 405792 18630
rect 405740 18566 405792 18572
rect 405844 16574 405872 18702
rect 405844 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 14482 407160 326402
rect 407212 326324 407264 326330
rect 407212 326266 407264 326272
rect 407224 225622 407252 326266
rect 407316 294642 407344 338014
rect 407592 326466 407620 338014
rect 407580 326460 407632 326466
rect 407580 326402 407632 326408
rect 407960 326330 407988 338014
rect 408558 337770 408586 338028
rect 408696 338014 408940 338042
rect 409064 338014 409308 338042
rect 409432 338014 409676 338042
rect 408558 337742 408632 337770
rect 408604 333198 408632 337742
rect 408592 333192 408644 333198
rect 408592 333134 408644 333140
rect 408696 330562 408724 338014
rect 408500 330540 408552 330546
rect 408500 330482 408552 330488
rect 408604 330534 408724 330562
rect 409064 330546 409092 338014
rect 409052 330540 409104 330546
rect 407948 326324 408000 326330
rect 407948 326266 408000 326272
rect 407304 294636 407356 294642
rect 407304 294578 407356 294584
rect 407212 225616 407264 225622
rect 407212 225558 407264 225564
rect 408512 25566 408540 330482
rect 408604 291854 408632 330534
rect 409052 330482 409104 330488
rect 409432 316034 409460 338014
rect 410030 337770 410058 338028
rect 410398 337770 410426 338028
rect 410536 338014 410780 338042
rect 410904 338014 411148 338042
rect 411272 338014 411516 338042
rect 411824 338014 411884 338042
rect 412008 338014 412252 338042
rect 412376 338014 412620 338042
rect 412744 338014 412988 338042
rect 413112 338014 413356 338042
rect 413480 338014 413724 338042
rect 410030 337742 410104 337770
rect 410398 337742 410472 337770
rect 409972 330540 410024 330546
rect 409972 330482 410024 330488
rect 408696 316006 409460 316034
rect 408696 308446 408724 316006
rect 408684 308440 408736 308446
rect 408684 308382 408736 308388
rect 409880 298784 409932 298790
rect 409880 298726 409932 298732
rect 408592 291848 408644 291854
rect 408592 291790 408644 291796
rect 408592 283688 408644 283694
rect 408592 283630 408644 283636
rect 407212 25560 407264 25566
rect 407212 25502 407264 25508
rect 408500 25560 408552 25566
rect 408500 25502 408552 25508
rect 407120 14476 407172 14482
rect 407120 14418 407172 14424
rect 407224 480 407252 25502
rect 408604 16574 408632 283630
rect 409892 16574 409920 298726
rect 409984 249082 410012 330482
rect 410076 290494 410104 337742
rect 410444 330478 410472 337742
rect 410432 330472 410484 330478
rect 410432 330414 410484 330420
rect 410536 316034 410564 338014
rect 410904 330546 410932 338014
rect 410892 330540 410944 330546
rect 410892 330482 410944 330488
rect 410168 316006 410564 316034
rect 410168 293282 410196 316006
rect 410156 293276 410208 293282
rect 410156 293218 410208 293224
rect 410064 290488 410116 290494
rect 410064 290430 410116 290436
rect 409972 249076 410024 249082
rect 409972 249018 410024 249024
rect 411272 32434 411300 338014
rect 411824 335510 411852 338014
rect 411812 335504 411864 335510
rect 411812 335446 411864 335452
rect 411352 330540 411404 330546
rect 411352 330482 411404 330488
rect 411364 224262 411392 330482
rect 412008 316034 412036 338014
rect 412376 330546 412404 338014
rect 412744 336682 412772 338014
rect 412652 336654 412772 336682
rect 412364 330540 412416 330546
rect 412364 330482 412416 330488
rect 411456 316006 412036 316034
rect 411456 289134 411484 316006
rect 411444 289128 411496 289134
rect 411444 289070 411496 289076
rect 411352 224256 411404 224262
rect 411352 224198 411404 224204
rect 411260 32428 411312 32434
rect 411260 32370 411312 32376
rect 408604 16546 409184 16574
rect 409892 16546 410840 16574
rect 408408 3596 408460 3602
rect 408408 3538 408460 3544
rect 408420 480 408448 3538
rect 404790 354 404902 480
rect 404464 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 412652 6186 412680 336654
rect 413112 335354 413140 338014
rect 413480 336682 413508 338014
rect 414078 337770 414106 338028
rect 414216 338014 414460 338042
rect 414584 338014 414828 338042
rect 414078 337742 414152 337770
rect 412744 335326 413140 335354
rect 413204 336654 413508 336682
rect 412744 8974 412772 335326
rect 413204 316034 413232 336654
rect 413284 335504 413336 335510
rect 413284 335446 413336 335452
rect 412836 316006 413232 316034
rect 412836 278050 412864 316006
rect 413296 304298 413324 335446
rect 413284 304292 413336 304298
rect 413284 304234 413336 304240
rect 412824 278044 412876 278050
rect 412824 277986 412876 277992
rect 412824 17264 412876 17270
rect 412824 17206 412876 17212
rect 412732 8968 412784 8974
rect 412732 8910 412784 8916
rect 412640 6180 412692 6186
rect 412640 6122 412692 6128
rect 411904 3460 411956 3466
rect 411904 3402 411956 3408
rect 411916 480 411944 3402
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412836 354 412864 17206
rect 414020 11756 414072 11762
rect 414020 11698 414072 11704
rect 414032 3074 414060 11698
rect 414124 3194 414152 337742
rect 414216 3602 414244 338014
rect 414584 316034 414612 338014
rect 414308 316006 414612 316034
rect 414308 16574 414336 316006
rect 414952 20670 414980 457422
rect 415400 282260 415452 282266
rect 415400 282202 415452 282208
rect 414940 20664 414992 20670
rect 414940 20606 414992 20612
rect 414308 16546 414428 16574
rect 414204 3596 414256 3602
rect 414204 3538 414256 3544
rect 414400 3369 414428 16546
rect 415412 3466 415440 282202
rect 417436 46918 417464 458322
rect 417528 431934 417556 461246
rect 422944 461236 422996 461242
rect 422944 461178 422996 461184
rect 421564 461168 421616 461174
rect 421564 461110 421616 461116
rect 420184 458516 420236 458522
rect 420184 458458 420236 458464
rect 418804 458448 418856 458454
rect 418804 458390 418856 458396
rect 417516 431928 417568 431934
rect 417516 431870 417568 431876
rect 417516 336456 417568 336462
rect 417516 336398 417568 336404
rect 417424 46912 417476 46918
rect 417424 46854 417476 46860
rect 416780 46232 416832 46238
rect 416780 46174 416832 46180
rect 416792 16574 416820 46174
rect 416792 16546 417464 16574
rect 415492 13116 415544 13122
rect 415492 13058 415544 13064
rect 415400 3460 415452 3466
rect 415400 3402 415452 3408
rect 414386 3360 414442 3369
rect 414386 3295 414442 3304
rect 414112 3188 414164 3194
rect 414112 3130 414164 3136
rect 414032 3046 414336 3074
rect 414308 480 414336 3046
rect 415504 480 415532 13058
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 416780 3460 416832 3466
rect 416780 3402 416832 3408
rect 416700 480 416728 3402
rect 416792 3194 416820 3402
rect 416780 3188 416832 3194
rect 416780 3130 416832 3136
rect 413070 354 413182 480
rect 412836 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417528 13122 417556 336398
rect 418816 86970 418844 458390
rect 419540 326392 419592 326398
rect 419540 326334 419592 326340
rect 418804 86964 418856 86970
rect 418804 86906 418856 86912
rect 419552 16574 419580 326334
rect 420196 167006 420224 458458
rect 421576 353258 421604 461110
rect 422956 405686 422984 461178
rect 424324 458720 424376 458726
rect 424324 458662 424376 458668
rect 422944 405680 422996 405686
rect 422944 405622 422996 405628
rect 424336 379506 424364 458662
rect 424324 379500 424376 379506
rect 424324 379442 424376 379448
rect 425716 365702 425744 462402
rect 462332 460766 462360 703520
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 478144 700324 478196 700330
rect 478144 700266 478196 700272
rect 478156 461650 478184 700266
rect 494072 464370 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 464364 494112 464370
rect 494060 464306 494112 464312
rect 478144 461644 478196 461650
rect 478144 461586 478196 461592
rect 462320 460760 462372 460766
rect 462320 460702 462372 460708
rect 527192 460630 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 460624 527232 460630
rect 527180 460566 527232 460572
rect 542372 460562 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 542360 460556 542412 460562
rect 542360 460498 542412 460504
rect 580264 458312 580316 458318
rect 580264 458254 580316 458260
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 427084 456884 427136 456890
rect 427084 456826 427136 456832
rect 427096 419490 427124 456826
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 427084 419484 427136 419490
rect 427084 419426 427136 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 425704 365696 425756 365702
rect 425704 365638 425756 365644
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 421564 353252 421616 353258
rect 421564 353194 421616 353200
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 424324 336388 424376 336394
rect 424324 336330 424376 336336
rect 421562 330440 421618 330449
rect 421562 330375 421618 330384
rect 420920 258732 420972 258738
rect 420920 258674 420972 258680
rect 420184 167000 420236 167006
rect 420184 166942 420236 166948
rect 419552 16546 420224 16574
rect 417516 13116 417568 13122
rect 417516 13058 417568 13064
rect 418988 3256 419040 3262
rect 418988 3198 419040 3204
rect 419000 480 419028 3198
rect 420196 480 420224 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 258674
rect 421576 206990 421604 330375
rect 422942 329080 422998 329089
rect 422942 329015 422998 329024
rect 422956 245614 422984 329015
rect 423680 324964 423732 324970
rect 423680 324906 423732 324912
rect 422944 245608 422996 245614
rect 422944 245550 422996 245556
rect 421564 206984 421616 206990
rect 421564 206926 421616 206932
rect 422576 3324 422628 3330
rect 422576 3266 422628 3272
rect 422588 480 422616 3266
rect 423692 1018 423720 324906
rect 423772 280900 423824 280906
rect 423772 280842 423824 280848
rect 423680 1012 423732 1018
rect 423680 954 423732 960
rect 423784 480 423812 280842
rect 424336 11762 424364 336330
rect 447140 336320 447192 336326
rect 447140 336262 447192 336268
rect 435362 331800 435418 331809
rect 435362 331735 435418 331744
rect 424414 327720 424470 327729
rect 424414 327655 424470 327664
rect 424428 299470 424456 327655
rect 425702 323640 425758 323649
rect 425702 323575 425758 323584
rect 424416 299464 424468 299470
rect 424416 299406 424468 299412
rect 425716 73166 425744 323575
rect 427082 322144 427138 322153
rect 427082 322079 427138 322088
rect 426440 279540 426492 279546
rect 426440 279482 426492 279488
rect 425704 73160 425756 73166
rect 425704 73102 425756 73108
rect 426452 16574 426480 279482
rect 427096 113150 427124 322079
rect 427820 320952 427872 320958
rect 427820 320894 427872 320900
rect 427084 113144 427136 113150
rect 427084 113086 427136 113092
rect 427832 16574 427860 320894
rect 434720 319524 434772 319530
rect 434720 319466 434772 319472
rect 428462 309768 428518 309777
rect 428462 309703 428518 309712
rect 428476 153202 428504 309703
rect 429842 308408 429898 308417
rect 429842 308343 429898 308352
rect 429856 193186 429884 308343
rect 431222 304192 431278 304201
rect 431222 304127 431278 304136
rect 431236 273222 431264 304127
rect 432602 301472 432658 301481
rect 432602 301407 432658 301416
rect 431224 273216 431276 273222
rect 431224 273158 431276 273164
rect 432052 247716 432104 247722
rect 432052 247658 432104 247664
rect 429844 193180 429896 193186
rect 429844 193122 429896 193128
rect 428464 153196 428516 153202
rect 428464 153138 428516 153144
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 424324 11756 424376 11762
rect 424324 11698 424376 11704
rect 426164 3392 426216 3398
rect 426164 3334 426216 3340
rect 424968 1012 425020 1018
rect 424968 954 425020 960
rect 424980 480 425008 954
rect 426176 480 426204 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 430856 6520 430908 6526
rect 430856 6462 430908 6468
rect 429660 4140 429712 4146
rect 429660 4082 429712 4088
rect 429672 480 429700 4082
rect 430868 480 430896 6462
rect 432064 480 432092 247658
rect 432616 60722 432644 301407
rect 432604 60716 432656 60722
rect 432604 60658 432656 60664
rect 434732 16574 434760 319466
rect 435376 126954 435404 331735
rect 441620 318164 441672 318170
rect 441620 318106 441672 318112
rect 438860 312588 438912 312594
rect 438860 312530 438912 312536
rect 438122 307048 438178 307057
rect 438122 306983 438178 306992
rect 436742 300112 436798 300121
rect 436742 300047 436798 300056
rect 435364 126948 435416 126954
rect 435364 126890 435416 126896
rect 436756 100706 436784 300047
rect 438136 233238 438164 306983
rect 438124 233232 438176 233238
rect 438124 233174 438176 233180
rect 436744 100700 436796 100706
rect 436744 100642 436796 100648
rect 438872 16574 438900 312530
rect 439502 291816 439558 291825
rect 439502 291751 439558 291760
rect 439516 139398 439544 291751
rect 440882 290456 440938 290465
rect 440882 290391 440938 290400
rect 440896 179382 440924 290391
rect 440884 179376 440936 179382
rect 440884 179318 440936 179324
rect 439504 139392 439556 139398
rect 439504 139334 439556 139340
rect 441632 16574 441660 318106
rect 442262 289096 442318 289105
rect 442262 289031 442318 289040
rect 442276 219434 442304 289031
rect 443642 287736 443698 287745
rect 443642 287671 443698 287680
rect 443656 259418 443684 287671
rect 443644 259412 443696 259418
rect 443644 259354 443696 259360
rect 442264 219428 442316 219434
rect 442264 219370 442316 219376
rect 447152 16574 447180 336262
rect 454040 336252 454092 336258
rect 454040 336194 454092 336200
rect 448520 278112 448572 278118
rect 448520 278054 448572 278060
rect 434732 16546 435128 16574
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 447152 16546 447456 16574
rect 434444 6452 434496 6458
rect 434444 6394 434496 6400
rect 433248 4072 433300 4078
rect 433248 4014 433300 4020
rect 433260 480 433288 4014
rect 434456 480 434484 6394
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 437940 6384 437992 6390
rect 437940 6326 437992 6332
rect 436744 4004 436796 4010
rect 436744 3946 436796 3952
rect 436756 480 436784 3946
rect 437952 480 437980 6326
rect 439148 480 439176 16546
rect 441528 6316 441580 6322
rect 441528 6258 441580 6264
rect 440332 3936 440384 3942
rect 440332 3878 440384 3884
rect 440344 480 440372 3878
rect 441540 480 441568 6258
rect 442644 480 442672 16546
rect 445760 10872 445812 10878
rect 445760 10814 445812 10820
rect 445024 6248 445076 6254
rect 445024 6190 445076 6196
rect 443828 3868 443880 3874
rect 443828 3810 443880 3816
rect 443840 480 443868 3810
rect 445036 480 445064 6190
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 10814
rect 447428 480 447456 16546
rect 448532 3210 448560 278054
rect 451280 276684 451332 276690
rect 451280 276626 451332 276632
rect 451292 16574 451320 276626
rect 451292 16546 451688 16574
rect 448612 10804 448664 10810
rect 448612 10746 448664 10752
rect 448624 3398 448652 10746
rect 450912 3800 450964 3806
rect 450912 3742 450964 3748
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 3742
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453304 10736 453356 10742
rect 453304 10678 453356 10684
rect 453316 480 453344 10678
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 336194
rect 460940 336184 460992 336190
rect 460940 336126 460992 336132
rect 455420 275324 455472 275330
rect 455420 275266 455472 275272
rect 455432 16574 455460 275266
rect 458180 273964 458232 273970
rect 458180 273906 458232 273912
rect 458192 16574 458220 273906
rect 460952 16574 460980 336126
rect 467840 336116 467892 336122
rect 467840 336058 467892 336064
rect 462320 286340 462372 286346
rect 462320 286282 462372 286288
rect 455432 16546 455736 16574
rect 458192 16546 459232 16574
rect 460952 16546 461624 16574
rect 455708 480 455736 16546
rect 456892 10668 456944 10674
rect 456892 10610 456944 10616
rect 456904 480 456932 10610
rect 458088 3732 458140 3738
rect 458088 3674 458140 3680
rect 458100 480 458128 3674
rect 459204 480 459232 16546
rect 459928 10600 459980 10606
rect 459928 10542 459980 10548
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 10542
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 286282
rect 465172 284980 465224 284986
rect 465172 284922 465224 284928
rect 465184 16574 465212 284922
rect 467852 16574 467880 336058
rect 474740 336048 474792 336054
rect 474740 335990 474792 335996
rect 473360 307080 473412 307086
rect 473360 307022 473412 307028
rect 470600 305720 470652 305726
rect 470600 305662 470652 305668
rect 469220 271176 469272 271182
rect 469220 271118 469272 271124
rect 469232 16574 469260 271118
rect 465184 16546 465856 16574
rect 467852 16546 468248 16574
rect 469232 16546 469904 16574
rect 463976 10532 464028 10538
rect 463976 10474 464028 10480
rect 463988 480 464016 10474
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 465184 480 465212 3606
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467472 10464 467524 10470
rect 467472 10406 467524 10412
rect 467484 480 467512 10406
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469876 480 469904 16546
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 305662
rect 473372 16574 473400 307022
rect 474752 16574 474780 335990
rect 480260 334688 480312 334694
rect 480260 334630 480312 334636
rect 480272 16574 480300 334630
rect 550640 334620 550692 334626
rect 550640 334562 550692 334568
rect 483020 333328 483072 333334
rect 483020 333270 483072 333276
rect 481640 269816 481692 269822
rect 481640 269758 481692 269764
rect 473372 16546 473492 16574
rect 474752 16546 475792 16574
rect 480272 16546 480576 16574
rect 472256 3528 472308 3534
rect 472256 3470 472308 3476
rect 472268 480 472296 3470
rect 473464 480 473492 16546
rect 474096 10396 474148 10402
rect 474096 10338 474148 10344
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 10338
rect 475764 480 475792 16546
rect 478144 10328 478196 10334
rect 478144 10270 478196 10276
rect 476948 7608 477000 7614
rect 476948 7550 477000 7556
rect 476960 480 476988 7550
rect 478156 480 478184 10270
rect 479338 3496 479394 3505
rect 479338 3431 479394 3440
rect 479352 480 479380 3431
rect 480548 480 480576 16546
rect 481652 6914 481680 269758
rect 481732 21412 481784 21418
rect 481732 21354 481784 21360
rect 481744 16574 481772 21354
rect 483032 16574 483060 333270
rect 525800 331900 525852 331906
rect 525800 331842 525852 331848
rect 500960 330608 501012 330614
rect 500960 330550 501012 330556
rect 487160 320884 487212 320890
rect 487160 320826 487212 320832
rect 484400 268388 484452 268394
rect 484400 268330 484452 268336
rect 484412 16574 484440 268330
rect 485780 246356 485832 246362
rect 485780 246298 485832 246304
rect 485792 16574 485820 246298
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 320826
rect 489920 319456 489972 319462
rect 489920 319398 489972 319404
rect 488540 267028 488592 267034
rect 488540 266970 488592 266976
rect 488552 16574 488580 266970
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 3534 489960 319398
rect 494060 318096 494112 318102
rect 494060 318038 494112 318044
rect 491300 265668 491352 265674
rect 491300 265610 491352 265616
rect 490012 24132 490064 24138
rect 490012 24074 490064 24080
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 24074
rect 491312 16574 491340 265610
rect 492680 243568 492732 243574
rect 492680 243510 492732 243516
rect 492692 16574 492720 243510
rect 494072 16574 494100 318038
rect 498200 316736 498252 316742
rect 498200 316678 498252 316684
rect 495440 264240 495492 264246
rect 495440 264182 495492 264188
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 264182
rect 496820 242208 496872 242214
rect 496820 242150 496872 242156
rect 496832 16574 496860 242150
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 316678
rect 498292 262880 498344 262886
rect 498292 262822 498344 262828
rect 498304 16574 498332 262822
rect 499580 240780 499632 240786
rect 499580 240722 499632 240728
rect 499592 16574 499620 240722
rect 500972 16574 501000 330550
rect 507860 329112 507912 329118
rect 507860 329054 507912 329060
rect 505100 305652 505152 305658
rect 505100 305594 505152 305600
rect 502340 261520 502392 261526
rect 502340 261462 502392 261468
rect 502352 16574 502380 261462
rect 503720 239420 503772 239426
rect 503720 239362 503772 239368
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 239362
rect 505112 16574 505140 305594
rect 506480 283620 506532 283626
rect 506480 283562 506532 283568
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 283562
rect 506572 26920 506624 26926
rect 506572 26862 506624 26868
rect 506584 16574 506612 26862
rect 507872 16574 507900 329054
rect 514760 327752 514812 327758
rect 514760 327694 514812 327700
rect 512000 313948 512052 313954
rect 512000 313890 512052 313896
rect 509240 260160 509292 260166
rect 509240 260102 509292 260108
rect 509252 16574 509280 260102
rect 510620 238060 510672 238066
rect 510620 238002 510672 238008
rect 510632 16574 510660 238002
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 313890
rect 513380 301504 513432 301510
rect 513380 301446 513432 301452
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 301446
rect 514772 3534 514800 327694
rect 518900 315308 518952 315314
rect 518900 315250 518952 315256
rect 516140 257372 516192 257378
rect 516140 257314 516192 257320
rect 514852 28280 514904 28286
rect 514852 28222 514904 28228
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 28222
rect 516152 16574 516180 257314
rect 517520 236700 517572 236706
rect 517520 236642 517572 236648
rect 517532 16574 517560 236642
rect 518912 16574 518940 315250
rect 520280 282192 520332 282198
rect 520280 282134 520332 282140
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 282134
rect 521660 235272 521712 235278
rect 521660 235214 521712 235220
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 235214
rect 524420 233912 524472 233918
rect 524420 233854 524472 233860
rect 523040 51740 523092 51746
rect 523040 51682 523092 51688
rect 523052 3534 523080 51682
rect 524432 16574 524460 233854
rect 525812 16574 525840 331842
rect 529940 323604 529992 323610
rect 529940 323546 529992 323552
rect 527180 300144 527232 300150
rect 527180 300086 527232 300092
rect 527192 16574 527220 300086
rect 528560 287700 528612 287706
rect 528560 287642 528612 287648
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523132 11756 523184 11762
rect 523132 11698 523184 11704
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 11698
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 287642
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 323546
rect 532700 322244 532752 322250
rect 532700 322186 532752 322192
rect 531320 256012 531372 256018
rect 531320 255954 531372 255960
rect 531332 480 531360 255954
rect 531412 22772 531464 22778
rect 531412 22714 531464 22720
rect 531424 16574 531452 22714
rect 532712 16574 532740 322186
rect 536840 311160 536892 311166
rect 536840 311102 536892 311108
rect 534080 254584 534132 254590
rect 534080 254526 534132 254532
rect 534092 16574 534120 254526
rect 535460 29640 535512 29646
rect 535460 29582 535512 29588
rect 535472 16574 535500 29582
rect 536852 16574 536880 311102
rect 543740 297424 543792 297430
rect 543740 297366 543792 297372
rect 538220 253224 538272 253230
rect 538220 253166 538272 253172
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 253166
rect 539600 231124 539652 231130
rect 539600 231066 539652 231072
rect 539612 480 539640 231066
rect 542360 229764 542412 229770
rect 542360 229706 542412 229712
rect 542372 16574 542400 229706
rect 543752 16574 543780 297366
rect 547880 295996 547932 296002
rect 547880 295938 547932 295944
rect 545120 251864 545172 251870
rect 545120 251806 545172 251812
rect 545132 16574 545160 251806
rect 546500 228404 546552 228410
rect 546500 228346 546552 228352
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 541992 13116 542044 13122
rect 541992 13058 542044 13064
rect 540796 4820 540848 4826
rect 540796 4762 540848 4768
rect 540808 480 540836 4762
rect 542004 480 542032 13058
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 228346
rect 547892 480 547920 295938
rect 547972 250504 548024 250510
rect 547972 250446 548024 250452
rect 547984 16574 548012 250446
rect 550652 16574 550680 334562
rect 561680 333260 561732 333266
rect 561680 333202 561732 333208
rect 554780 309800 554832 309806
rect 554780 309742 554832 309748
rect 552020 280832 552072 280838
rect 552020 280774 552072 280780
rect 552032 16574 552060 280774
rect 553400 227044 553452 227050
rect 553400 226986 553452 226992
rect 553412 16574 553440 226986
rect 547984 16546 548656 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550272 15904 550324 15910
rect 550272 15846 550324 15852
rect 550284 480 550312 15846
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 309742
rect 557540 294636 557592 294642
rect 557540 294578 557592 294584
rect 556160 279472 556212 279478
rect 556160 279414 556212 279420
rect 556172 480 556200 279414
rect 556252 18624 556304 18630
rect 556252 18566 556304 18572
rect 556264 16574 556292 18566
rect 557552 16574 557580 294578
rect 560300 225616 560352 225622
rect 560300 225558 560352 225564
rect 560312 16574 560340 225558
rect 561692 16574 561720 333202
rect 567200 330540 567252 330546
rect 567200 330482 567252 330488
rect 564440 308440 564492 308446
rect 564440 308382 564492 308388
rect 563060 291848 563112 291854
rect 563060 291790 563112 291796
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 559288 14476 559340 14482
rect 559288 14418 559340 14424
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 14418
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 291790
rect 564452 3534 564480 308382
rect 565820 290488 565872 290494
rect 565820 290430 565872 290436
rect 564532 25560 564584 25566
rect 564532 25502 564584 25508
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 25502
rect 565832 16574 565860 290430
rect 567212 16574 567240 330482
rect 572812 304292 572864 304298
rect 572812 304234 572864 304240
rect 568580 293276 568632 293282
rect 568580 293218 568632 293224
rect 568592 16574 568620 293218
rect 571984 289128 572036 289134
rect 571984 289070 572036 289076
rect 569960 249076 570012 249082
rect 569960 249018 570012 249024
rect 569972 16574 570000 249018
rect 571340 32428 571392 32434
rect 571340 32370 571392 32376
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 32370
rect 571996 3058 572024 289070
rect 572824 6914 572852 304234
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 576124 278044 576176 278050
rect 576124 277986 576176 277992
rect 574100 224256 574152 224262
rect 574100 224198 574152 224204
rect 574112 16574 574140 224198
rect 574112 16546 575152 16574
rect 572732 6886 572852 6914
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 6886
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 16546
rect 576136 3806 576164 277986
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 579712 100700 579764 100706
rect 579712 100642 579764 100648
rect 579724 99521 579752 100642
rect 579710 99512 579766 99521
rect 579710 99447 579766 99456
rect 579988 86964 580040 86970
rect 579988 86906 580040 86912
rect 580000 86193 580028 86906
rect 579986 86184 580042 86193
rect 579986 86119 580042 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 579804 60716 579856 60722
rect 579804 60658 579856 60664
rect 579816 59673 579844 60658
rect 579802 59664 579858 59673
rect 579802 59599 579858 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576124 3800 576176 3806
rect 576124 3742 576176 3748
rect 576320 480 576348 6122
rect 577424 480 577452 8910
rect 580276 6633 580304 458254
rect 580354 326360 580410 326369
rect 580354 326295 580410 326304
rect 580368 33153 580396 326295
rect 580446 302832 580502 302841
rect 580446 302767 580502 302776
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 580460 19825 580488 302767
rect 580446 19816 580502 19825
rect 580446 19751 580502 19760
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 578608 3800 578660 3806
rect 578608 3742 578660 3748
rect 578620 480 578648 3742
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 619112 3386 619168
rect 3330 606056 3386 606112
rect 3054 566888 3110 566944
rect 3330 553832 3386 553888
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632032 3570 632088
rect 3606 579944 3662 580000
rect 3698 527856 3754 527912
rect 3882 475632 3938 475688
rect 3514 462576 3570 462632
rect 3422 460128 3478 460184
rect 3330 449520 3386 449576
rect 2962 410488 3018 410544
rect 3606 423544 3662 423600
rect 3514 397432 3570 397488
rect 3514 371320 3570 371376
rect 3422 358400 3478 358456
rect 3146 345344 3202 345400
rect 3330 306176 3386 306232
rect 2870 293120 2926 293176
rect 3238 267144 3294 267200
rect 3330 254088 3386 254144
rect 3238 241032 3294 241088
rect 2778 214956 2780 214976
rect 2780 214956 2832 214976
rect 2832 214956 2834 214976
rect 2778 214920 2834 214956
rect 3330 201864 3386 201920
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3330 149776 3386 149832
rect 3238 110608 3294 110664
rect 3238 97552 3294 97608
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 3330 58520 3386 58576
rect 2778 32444 2780 32464
rect 2780 32444 2832 32464
rect 2832 32444 2834 32464
rect 2778 32408 2834 32444
rect 3514 319232 3570 319288
rect 3606 316648 3662 316704
rect 3514 313928 3570 313984
rect 3606 136720 3662 136776
rect 3514 45464 3570 45520
rect 3514 19352 3570 19408
rect 3514 6468 3516 6488
rect 3516 6468 3568 6488
rect 3568 6468 3570 6488
rect 3514 6432 3570 6468
rect 40038 460264 40094 460320
rect 7562 337320 7618 337376
rect 6182 333240 6238 333296
rect 5262 3304 5318 3360
rect 8942 311072 8998 311128
rect 11150 3440 11206 3496
rect 18602 320728 18658 320784
rect 11794 297336 11850 297392
rect 13174 295976 13230 296032
rect 14462 294480 14518 294536
rect 21362 315288 21418 315344
rect 40682 318008 40738 318064
rect 31022 298696 31078 298752
rect 28262 293120 28318 293176
rect 344374 460264 344430 460320
rect 349158 460128 349214 460184
rect 407578 459720 407634 459776
rect 237654 457408 237710 457464
rect 239218 457408 239274 457464
rect 242346 457408 242402 457464
rect 243910 457408 243966 457464
rect 246670 457408 246726 457464
rect 248234 457408 248290 457464
rect 250258 457408 250314 457464
rect 251822 457408 251878 457464
rect 253386 457408 253442 457464
rect 256514 457408 256570 457464
rect 257710 457408 257766 457464
rect 259274 457408 259330 457464
rect 261298 457408 261354 457464
rect 262862 457408 262918 457464
rect 264518 457408 264574 457464
rect 266082 457408 266138 457464
rect 267554 457408 267610 457464
rect 268750 457408 268806 457464
rect 270590 457408 270646 457464
rect 272338 457408 272394 457464
rect 383842 457408 383898 457464
rect 385406 457408 385462 457464
rect 388626 457408 388682 457464
rect 390190 457408 390246 457464
rect 393502 457408 393558 457464
rect 394882 457408 394938 457464
rect 398102 457408 398158 457464
rect 399666 457408 399722 457464
rect 401230 457408 401286 457464
rect 402978 457408 403034 457464
rect 404358 457408 404414 457464
rect 406014 457408 406070 457464
rect 409142 457408 409198 457464
rect 410706 457408 410762 457464
rect 412270 457408 412326 457464
rect 233882 334600 233938 334656
rect 232594 319368 232650 319424
rect 236274 3304 236330 3360
rect 237378 3440 237434 3496
rect 277122 3304 277178 3360
rect 320270 3304 320326 3360
rect 383014 336776 383070 336832
rect 382554 3440 382610 3496
rect 414386 3304 414442 3360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 579618 404912 579674 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 421562 330384 421618 330440
rect 422942 329024 422998 329080
rect 435362 331744 435418 331800
rect 424414 327664 424470 327720
rect 425702 323584 425758 323640
rect 427082 322088 427138 322144
rect 428462 309712 428518 309768
rect 429842 308352 429898 308408
rect 431222 304136 431278 304192
rect 432602 301416 432658 301472
rect 438122 306992 438178 307048
rect 436742 300056 436798 300112
rect 439502 291760 439558 291816
rect 440882 290400 440938 290456
rect 442262 289040 442318 289096
rect 443642 287680 443698 287736
rect 479338 3440 479394 3496
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579618 125976 579674 126032
rect 580170 112784 580226 112840
rect 579710 99456 579766 99512
rect 579986 86128 580042 86184
rect 580170 72936 580226 72992
rect 579802 59608 579858 59664
rect 580170 46280 580226 46336
rect 580354 326304 580410 326360
rect 580446 302776 580502 302832
rect 580354 33088 580410 33144
rect 580446 19760 580502 19816
rect 580262 6568 580318 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3325 619170 3391 619173
rect -960 619168 3391 619170
rect -960 619112 3330 619168
rect 3386 619112 3391 619168
rect -960 619110 3391 619112
rect -960 619020 480 619110
rect 3325 619107 3391 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3601 580002 3667 580005
rect -960 580000 3667 580002
rect -960 579944 3606 580000
rect 3662 579944 3667 580000
rect -960 579942 3667 579944
rect -960 579852 480 579942
rect 3601 579939 3667 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3693 527914 3759 527917
rect -960 527912 3759 527914
rect -960 527856 3698 527912
rect 3754 527856 3759 527912
rect -960 527854 3759 527856
rect -960 527764 480 527854
rect 3693 527851 3759 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 40033 460322 40099 460325
rect 344369 460322 344435 460325
rect 40033 460320 344435 460322
rect 40033 460264 40038 460320
rect 40094 460264 344374 460320
rect 344430 460264 344435 460320
rect 40033 460262 344435 460264
rect 40033 460259 40099 460262
rect 344369 460259 344435 460262
rect 3417 460186 3483 460189
rect 349153 460186 349219 460189
rect 3417 460184 349219 460186
rect 3417 460128 3422 460184
rect 3478 460128 349158 460184
rect 349214 460128 349219 460184
rect 3417 460126 349219 460128
rect 3417 460123 3483 460126
rect 349153 460123 349219 460126
rect 402094 459716 402100 459780
rect 402164 459778 402170 459780
rect 407573 459778 407639 459781
rect 402164 459776 407639 459778
rect 402164 459720 407578 459776
rect 407634 459720 407639 459776
rect 402164 459718 407639 459720
rect 402164 459716 402170 459718
rect 407573 459715 407639 459718
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 237649 457466 237715 457469
rect 237966 457466 237972 457468
rect 237649 457464 237972 457466
rect 237649 457408 237654 457464
rect 237710 457408 237972 457464
rect 237649 457406 237972 457408
rect 237649 457403 237715 457406
rect 237966 457404 237972 457406
rect 238036 457404 238042 457468
rect 239213 457466 239279 457469
rect 240726 457466 240732 457468
rect 239213 457464 240732 457466
rect 239213 457408 239218 457464
rect 239274 457408 240732 457464
rect 239213 457406 240732 457408
rect 239213 457403 239279 457406
rect 240726 457404 240732 457406
rect 240796 457404 240802 457468
rect 242341 457466 242407 457469
rect 242750 457466 242756 457468
rect 242341 457464 242756 457466
rect 242341 457408 242346 457464
rect 242402 457408 242756 457464
rect 242341 457406 242756 457408
rect 242341 457403 242407 457406
rect 242750 457404 242756 457406
rect 242820 457404 242826 457468
rect 243905 457466 243971 457469
rect 244038 457466 244044 457468
rect 243905 457464 244044 457466
rect 243905 457408 243910 457464
rect 243966 457408 244044 457464
rect 243905 457406 244044 457408
rect 243905 457403 243971 457406
rect 244038 457404 244044 457406
rect 244108 457404 244114 457468
rect 246665 457466 246731 457469
rect 248229 457468 248295 457469
rect 246798 457466 246804 457468
rect 246665 457464 246804 457466
rect 246665 457408 246670 457464
rect 246726 457408 246804 457464
rect 246665 457406 246804 457408
rect 246665 457403 246731 457406
rect 246798 457404 246804 457406
rect 246868 457404 246874 457468
rect 248229 457464 248276 457468
rect 248340 457466 248346 457468
rect 250253 457466 250319 457469
rect 251030 457466 251036 457468
rect 248229 457408 248234 457464
rect 248229 457404 248276 457408
rect 248340 457406 248386 457466
rect 250253 457464 251036 457466
rect 250253 457408 250258 457464
rect 250314 457408 251036 457464
rect 250253 457406 251036 457408
rect 248340 457404 248346 457406
rect 248229 457403 248295 457404
rect 250253 457403 250319 457406
rect 251030 457404 251036 457406
rect 251100 457404 251106 457468
rect 251817 457466 251883 457469
rect 252318 457466 252324 457468
rect 251817 457464 252324 457466
rect 251817 457408 251822 457464
rect 251878 457408 252324 457464
rect 251817 457406 252324 457408
rect 251817 457403 251883 457406
rect 252318 457404 252324 457406
rect 252388 457404 252394 457468
rect 253381 457466 253447 457469
rect 256509 457468 256575 457469
rect 253606 457466 253612 457468
rect 253381 457464 253612 457466
rect 253381 457408 253386 457464
rect 253442 457408 253612 457464
rect 253381 457406 253612 457408
rect 253381 457403 253447 457406
rect 253606 457404 253612 457406
rect 253676 457404 253682 457468
rect 256509 457464 256556 457468
rect 256620 457466 256626 457468
rect 257705 457466 257771 457469
rect 259269 457468 259335 457469
rect 257838 457466 257844 457468
rect 256509 457408 256514 457464
rect 256509 457404 256556 457408
rect 256620 457406 256666 457466
rect 257705 457464 257844 457466
rect 257705 457408 257710 457464
rect 257766 457408 257844 457464
rect 257705 457406 257844 457408
rect 256620 457404 256626 457406
rect 256509 457403 256575 457404
rect 257705 457403 257771 457406
rect 257838 457404 257844 457406
rect 257908 457404 257914 457468
rect 259269 457464 259316 457468
rect 259380 457466 259386 457468
rect 261293 457466 261359 457469
rect 262070 457466 262076 457468
rect 259269 457408 259274 457464
rect 259269 457404 259316 457408
rect 259380 457406 259426 457466
rect 261293 457464 262076 457466
rect 261293 457408 261298 457464
rect 261354 457408 262076 457464
rect 261293 457406 262076 457408
rect 259380 457404 259386 457406
rect 259269 457403 259335 457404
rect 261293 457403 261359 457406
rect 262070 457404 262076 457406
rect 262140 457404 262146 457468
rect 262857 457466 262923 457469
rect 263358 457466 263364 457468
rect 262857 457464 263364 457466
rect 262857 457408 262862 457464
rect 262918 457408 263364 457464
rect 262857 457406 263364 457408
rect 262857 457403 262923 457406
rect 263358 457404 263364 457406
rect 263428 457404 263434 457468
rect 264513 457466 264579 457469
rect 266077 457468 266143 457469
rect 267549 457468 267615 457469
rect 264830 457466 264836 457468
rect 264513 457464 264836 457466
rect 264513 457408 264518 457464
rect 264574 457408 264836 457464
rect 264513 457406 264836 457408
rect 264513 457403 264579 457406
rect 264830 457404 264836 457406
rect 264900 457404 264906 457468
rect 266077 457464 266124 457468
rect 266188 457466 266194 457468
rect 266077 457408 266082 457464
rect 266077 457404 266124 457408
rect 266188 457406 266234 457466
rect 267549 457464 267596 457468
rect 267660 457466 267666 457468
rect 268745 457466 268811 457469
rect 268878 457466 268884 457468
rect 267549 457408 267554 457464
rect 266188 457404 266194 457406
rect 267549 457404 267596 457408
rect 267660 457406 267706 457466
rect 268745 457464 268884 457466
rect 268745 457408 268750 457464
rect 268806 457408 268884 457464
rect 268745 457406 268884 457408
rect 267660 457404 267666 457406
rect 266077 457403 266143 457404
rect 267549 457403 267615 457404
rect 268745 457403 268811 457406
rect 268878 457404 268884 457406
rect 268948 457404 268954 457468
rect 270585 457466 270651 457469
rect 271086 457466 271092 457468
rect 270585 457464 271092 457466
rect 270585 457408 270590 457464
rect 270646 457408 271092 457464
rect 270585 457406 271092 457408
rect 270585 457403 270651 457406
rect 271086 457404 271092 457406
rect 271156 457404 271162 457468
rect 272333 457466 272399 457469
rect 273846 457466 273852 457468
rect 272333 457464 273852 457466
rect 272333 457408 272338 457464
rect 272394 457408 273852 457464
rect 272333 457406 273852 457408
rect 272333 457403 272399 457406
rect 273846 457404 273852 457406
rect 273916 457404 273922 457468
rect 383694 457404 383700 457468
rect 383764 457466 383770 457468
rect 383837 457466 383903 457469
rect 383764 457464 383903 457466
rect 383764 457408 383842 457464
rect 383898 457408 383903 457464
rect 383764 457406 383903 457408
rect 383764 457404 383770 457406
rect 383837 457403 383903 457406
rect 384982 457404 384988 457468
rect 385052 457466 385058 457468
rect 385401 457466 385467 457469
rect 385052 457464 385467 457466
rect 385052 457408 385406 457464
rect 385462 457408 385467 457464
rect 385052 457406 385467 457408
rect 385052 457404 385058 457406
rect 385401 457403 385467 457406
rect 387742 457404 387748 457468
rect 387812 457466 387818 457468
rect 388621 457466 388687 457469
rect 387812 457464 388687 457466
rect 387812 457408 388626 457464
rect 388682 457408 388687 457464
rect 387812 457406 388687 457408
rect 387812 457404 387818 457406
rect 388621 457403 388687 457406
rect 389214 457404 389220 457468
rect 389284 457466 389290 457468
rect 390185 457466 390251 457469
rect 393497 457468 393563 457469
rect 393446 457466 393452 457468
rect 389284 457464 390251 457466
rect 389284 457408 390190 457464
rect 390246 457408 390251 457464
rect 389284 457406 390251 457408
rect 393406 457406 393452 457466
rect 393516 457464 393563 457468
rect 393558 457408 393563 457464
rect 389284 457404 389290 457406
rect 390185 457403 390251 457406
rect 393446 457404 393452 457406
rect 393516 457404 393563 457408
rect 394734 457404 394740 457468
rect 394804 457466 394810 457468
rect 394877 457466 394943 457469
rect 394804 457464 394943 457466
rect 394804 457408 394882 457464
rect 394938 457408 394943 457464
rect 394804 457406 394943 457408
rect 394804 457404 394810 457406
rect 393497 457403 393563 457404
rect 394877 457403 394943 457406
rect 396574 457404 396580 457468
rect 396644 457466 396650 457468
rect 398097 457466 398163 457469
rect 396644 457464 398163 457466
rect 396644 457408 398102 457464
rect 398158 457408 398163 457464
rect 396644 457406 398163 457408
rect 396644 457404 396650 457406
rect 398097 457403 398163 457406
rect 398782 457404 398788 457468
rect 398852 457466 398858 457468
rect 399661 457466 399727 457469
rect 398852 457464 399727 457466
rect 398852 457408 399666 457464
rect 399722 457408 399727 457464
rect 398852 457406 399727 457408
rect 398852 457404 398858 457406
rect 399661 457403 399727 457406
rect 400254 457404 400260 457468
rect 400324 457466 400330 457468
rect 401225 457466 401291 457469
rect 400324 457464 401291 457466
rect 400324 457408 401230 457464
rect 401286 457408 401291 457464
rect 400324 457406 401291 457408
rect 400324 457404 400330 457406
rect 401225 457403 401291 457406
rect 402973 457468 403039 457469
rect 404353 457468 404419 457469
rect 402973 457464 403020 457468
rect 403084 457466 403090 457468
rect 404302 457466 404308 457468
rect 402973 457408 402978 457464
rect 402973 457404 403020 457408
rect 403084 457406 403130 457466
rect 404262 457406 404308 457466
rect 404372 457464 404419 457468
rect 404414 457408 404419 457464
rect 403084 457404 403090 457406
rect 404302 457404 404308 457406
rect 404372 457404 404419 457408
rect 405774 457404 405780 457468
rect 405844 457466 405850 457468
rect 406009 457466 406075 457469
rect 405844 457464 406075 457466
rect 405844 457408 406014 457464
rect 406070 457408 406075 457464
rect 405844 457406 406075 457408
rect 405844 457404 405850 457406
rect 402973 457403 403039 457404
rect 404353 457403 404419 457404
rect 406009 457403 406075 457406
rect 408718 457404 408724 457468
rect 408788 457466 408794 457468
rect 409137 457466 409203 457469
rect 408788 457464 409203 457466
rect 408788 457408 409142 457464
rect 409198 457408 409203 457464
rect 408788 457406 409203 457408
rect 408788 457404 408794 457406
rect 409137 457403 409203 457406
rect 409822 457404 409828 457468
rect 409892 457466 409898 457468
rect 410701 457466 410767 457469
rect 409892 457464 410767 457466
rect 409892 457408 410706 457464
rect 410762 457408 410767 457464
rect 409892 457406 410767 457408
rect 409892 457404 409898 457406
rect 410701 457403 410767 457406
rect 411294 457404 411300 457468
rect 411364 457466 411370 457468
rect 412265 457466 412331 457469
rect 411364 457464 412331 457466
rect 411364 457408 412270 457464
rect 412326 457408 412331 457464
rect 411364 457406 412331 457408
rect 411364 457404 411370 457406
rect 412265 457403 412331 457406
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3601 423602 3667 423605
rect -960 423600 3667 423602
rect -960 423544 3606 423600
rect 3662 423544 3667 423600
rect -960 423542 3667 423544
rect -960 423452 480 423542
rect 3601 423539 3667 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 583520 338452 584960 338692
rect 7557 337378 7623 337381
rect 400254 337378 400260 337380
rect 7557 337376 400260 337378
rect 7557 337320 7562 337376
rect 7618 337320 400260 337376
rect 7557 337318 400260 337320
rect 7557 337315 7623 337318
rect 400254 337316 400260 337318
rect 400324 337316 400330 337380
rect 383009 336834 383075 336837
rect 384982 336834 384988 336836
rect 383009 336832 384988 336834
rect 383009 336776 383014 336832
rect 383070 336776 384988 336832
rect 383009 336774 384988 336776
rect 383009 336771 383075 336774
rect 384982 336772 384988 336774
rect 385052 336772 385058 336836
rect 233877 334658 233943 334661
rect 405774 334658 405780 334660
rect 233877 334656 405780 334658
rect 233877 334600 233882 334656
rect 233938 334600 405780 334656
rect 233877 334598 405780 334600
rect 233877 334595 233943 334598
rect 405774 334596 405780 334598
rect 405844 334596 405850 334660
rect 6177 333298 6243 333301
rect 409822 333298 409828 333300
rect 6177 333296 409828 333298
rect 6177 333240 6182 333296
rect 6238 333240 409828 333296
rect 6177 333238 409828 333240
rect 6177 333235 6243 333238
rect 409822 333236 409828 333238
rect 409892 333236 409898 333300
rect -960 332196 480 332436
rect 251030 331740 251036 331804
rect 251100 331802 251106 331804
rect 435357 331802 435423 331805
rect 251100 331800 435423 331802
rect 251100 331744 435362 331800
rect 435418 331744 435423 331800
rect 251100 331742 435423 331744
rect 251100 331740 251106 331742
rect 435357 331739 435423 331742
rect 259310 330380 259316 330444
rect 259380 330442 259386 330444
rect 421557 330442 421623 330445
rect 259380 330440 421623 330442
rect 259380 330384 421562 330440
rect 421618 330384 421623 330440
rect 259380 330382 421623 330384
rect 259380 330380 259386 330382
rect 421557 330379 421623 330382
rect 264830 329020 264836 329084
rect 264900 329082 264906 329084
rect 422937 329082 423003 329085
rect 264900 329080 423003 329082
rect 264900 329024 422942 329080
rect 422998 329024 423003 329080
rect 264900 329022 423003 329024
rect 264900 329020 264906 329022
rect 422937 329019 423003 329022
rect 268878 327660 268884 327724
rect 268948 327722 268954 327724
rect 424409 327722 424475 327725
rect 268948 327720 424475 327722
rect 268948 327664 424414 327720
rect 424470 327664 424475 327720
rect 268948 327662 424475 327664
rect 268948 327660 268954 327662
rect 424409 327659 424475 327662
rect 237966 326300 237972 326364
rect 238036 326362 238042 326364
rect 580349 326362 580415 326365
rect 238036 326360 580415 326362
rect 238036 326304 580354 326360
rect 580410 326304 580415 326360
rect 238036 326302 580415 326304
rect 238036 326300 238042 326302
rect 580349 326299 580415 326302
rect 583520 325274 584960 325364
rect 583342 325214 584960 325274
rect 583342 325138 583402 325214
rect 583520 325138 584960 325214
rect 583342 325124 584960 325138
rect 583342 325078 583586 325124
rect 271086 324396 271092 324460
rect 271156 324458 271162 324460
rect 583526 324458 583586 325078
rect 271156 324398 583586 324458
rect 271156 324396 271162 324398
rect 242750 323580 242756 323644
rect 242820 323642 242826 323644
rect 425697 323642 425763 323645
rect 242820 323640 425763 323642
rect 242820 323584 425702 323640
rect 425758 323584 425763 323640
rect 242820 323582 425763 323584
rect 242820 323580 242826 323582
rect 425697 323579 425763 323582
rect 246798 322084 246804 322148
rect 246868 322146 246874 322148
rect 427077 322146 427143 322149
rect 246868 322144 427143 322146
rect 246868 322088 427082 322144
rect 427138 322088 427143 322144
rect 246868 322086 427143 322088
rect 246868 322084 246874 322086
rect 427077 322083 427143 322086
rect 18597 320786 18663 320789
rect 383694 320786 383700 320788
rect 18597 320784 383700 320786
rect 18597 320728 18602 320784
rect 18658 320728 383700 320784
rect 18597 320726 383700 320728
rect 18597 320723 18663 320726
rect 383694 320724 383700 320726
rect 383764 320724 383770 320788
rect 232589 319426 232655 319429
rect 387742 319426 387748 319428
rect 232589 319424 387748 319426
rect -960 319290 480 319380
rect 232589 319368 232594 319424
rect 232650 319368 387748 319424
rect 232589 319366 387748 319368
rect 232589 319363 232655 319366
rect 387742 319364 387748 319366
rect 387812 319364 387818 319428
rect 3509 319290 3575 319293
rect -960 319288 3575 319290
rect -960 319232 3514 319288
rect 3570 319232 3575 319288
rect -960 319230 3575 319232
rect -960 319140 480 319230
rect 3509 319227 3575 319230
rect 40677 318066 40743 318069
rect 393078 318066 393084 318068
rect 40677 318064 393084 318066
rect 40677 318008 40682 318064
rect 40738 318008 393084 318064
rect 40677 318006 393084 318008
rect 40677 318003 40743 318006
rect 393078 318004 393084 318006
rect 393148 318004 393154 318068
rect 3601 316706 3667 316709
rect 396574 316706 396580 316708
rect 3601 316704 396580 316706
rect 3601 316648 3606 316704
rect 3662 316648 396580 316704
rect 3601 316646 396580 316648
rect 3601 316643 3667 316646
rect 396574 316644 396580 316646
rect 396644 316644 396650 316708
rect 21357 315346 21423 315349
rect 403014 315346 403020 315348
rect 21357 315344 403020 315346
rect 21357 315288 21362 315344
rect 21418 315288 403020 315344
rect 21357 315286 403020 315288
rect 21357 315283 21423 315286
rect 403014 315284 403020 315286
rect 403084 315284 403090 315348
rect 3509 313986 3575 313989
rect 402094 313986 402100 313988
rect 3509 313984 402100 313986
rect 3509 313928 3514 313984
rect 3570 313928 402100 313984
rect 3509 313926 402100 313928
rect 3509 313923 3575 313926
rect 402094 313924 402100 313926
rect 402164 313924 402170 313988
rect 583520 312082 584960 312172
rect 567150 312022 584960 312082
rect 273846 311884 273852 311948
rect 273916 311946 273922 311948
rect 567150 311946 567210 312022
rect 273916 311886 567210 311946
rect 583520 311932 584960 312022
rect 273916 311884 273922 311886
rect 8937 311130 9003 311133
rect 411294 311130 411300 311132
rect 8937 311128 411300 311130
rect 8937 311072 8942 311128
rect 8998 311072 411300 311128
rect 8937 311070 411300 311072
rect 8937 311067 9003 311070
rect 411294 311068 411300 311070
rect 411364 311068 411370 311132
rect 252318 309708 252324 309772
rect 252388 309770 252394 309772
rect 428457 309770 428523 309773
rect 252388 309768 428523 309770
rect 252388 309712 428462 309768
rect 428518 309712 428523 309768
rect 252388 309710 428523 309712
rect 252388 309708 252394 309710
rect 428457 309707 428523 309710
rect 256550 308348 256556 308412
rect 256620 308410 256626 308412
rect 429837 308410 429903 308413
rect 256620 308408 429903 308410
rect 256620 308352 429842 308408
rect 429898 308352 429903 308408
rect 256620 308350 429903 308352
rect 256620 308348 256626 308350
rect 429837 308347 429903 308350
rect 262070 306988 262076 307052
rect 262140 307050 262146 307052
rect 438117 307050 438183 307053
rect 262140 307048 438183 307050
rect 262140 306992 438122 307048
rect 438178 306992 438183 307048
rect 262140 306990 438183 306992
rect 262140 306988 262146 306990
rect 438117 306987 438183 306990
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 266118 304132 266124 304196
rect 266188 304194 266194 304196
rect 431217 304194 431283 304197
rect 266188 304192 431283 304194
rect 266188 304136 431222 304192
rect 431278 304136 431283 304192
rect 266188 304134 431283 304136
rect 266188 304132 266194 304134
rect 431217 304131 431283 304134
rect 240726 302772 240732 302836
rect 240796 302834 240802 302836
rect 580441 302834 580507 302837
rect 240796 302832 580507 302834
rect 240796 302776 580446 302832
rect 580502 302776 580507 302832
rect 240796 302774 580507 302776
rect 240796 302772 240802 302774
rect 580441 302771 580507 302774
rect 244038 301412 244044 301476
rect 244108 301474 244114 301476
rect 432597 301474 432663 301477
rect 244108 301472 432663 301474
rect 244108 301416 432602 301472
rect 432658 301416 432663 301472
rect 244108 301414 432663 301416
rect 244108 301412 244114 301414
rect 432597 301411 432663 301414
rect 248270 300052 248276 300116
rect 248340 300114 248346 300116
rect 436737 300114 436803 300117
rect 248340 300112 436803 300114
rect 248340 300056 436742 300112
rect 436798 300056 436803 300112
rect 248340 300054 436803 300056
rect 248340 300052 248346 300054
rect 436737 300051 436803 300054
rect 31017 298754 31083 298757
rect 389214 298754 389220 298756
rect 31017 298752 389220 298754
rect 31017 298696 31022 298752
rect 31078 298696 389220 298752
rect 31017 298694 389220 298696
rect 31017 298691 31083 298694
rect 389214 298692 389220 298694
rect 389284 298692 389290 298756
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 11789 297394 11855 297397
rect 394734 297394 394740 297396
rect 11789 297392 394740 297394
rect 11789 297336 11794 297392
rect 11850 297336 394740 297392
rect 11789 297334 394740 297336
rect 11789 297331 11855 297334
rect 394734 297332 394740 297334
rect 394804 297332 394810 297396
rect 13169 296034 13235 296037
rect 398782 296034 398788 296036
rect 13169 296032 398788 296034
rect 13169 295976 13174 296032
rect 13230 295976 398788 296032
rect 13169 295974 398788 295976
rect 13169 295971 13235 295974
rect 398782 295972 398788 295974
rect 398852 295972 398858 296036
rect 14457 294538 14523 294541
rect 404302 294538 404308 294540
rect 14457 294536 404308 294538
rect 14457 294480 14462 294536
rect 14518 294480 404308 294536
rect 14457 294478 404308 294480
rect 14457 294475 14523 294478
rect 404302 294476 404308 294478
rect 404372 294476 404378 294540
rect -960 293178 480 293268
rect 2865 293178 2931 293181
rect -960 293176 2931 293178
rect -960 293120 2870 293176
rect 2926 293120 2931 293176
rect -960 293118 2931 293120
rect -960 293028 480 293118
rect 2865 293115 2931 293118
rect 28257 293178 28323 293181
rect 408718 293178 408724 293180
rect 28257 293176 408724 293178
rect 28257 293120 28262 293176
rect 28318 293120 408724 293176
rect 28257 293118 408724 293120
rect 28257 293115 28323 293118
rect 408718 293116 408724 293118
rect 408788 293116 408794 293180
rect 253606 291756 253612 291820
rect 253676 291818 253682 291820
rect 439497 291818 439563 291821
rect 253676 291816 439563 291818
rect 253676 291760 439502 291816
rect 439558 291760 439563 291816
rect 253676 291758 439563 291760
rect 253676 291756 253682 291758
rect 439497 291755 439563 291758
rect 257838 290396 257844 290460
rect 257908 290458 257914 290460
rect 440877 290458 440943 290461
rect 257908 290456 440943 290458
rect 257908 290400 440882 290456
rect 440938 290400 440943 290456
rect 257908 290398 440943 290400
rect 257908 290396 257914 290398
rect 440877 290395 440943 290398
rect 263358 289036 263364 289100
rect 263428 289098 263434 289100
rect 442257 289098 442323 289101
rect 263428 289096 442323 289098
rect 263428 289040 442262 289096
rect 442318 289040 442323 289096
rect 263428 289038 442323 289040
rect 263428 289036 263434 289038
rect 442257 289035 442323 289038
rect 267590 287676 267596 287740
rect 267660 287738 267666 287740
rect 443637 287738 443703 287741
rect 267660 287736 443703 287738
rect 267660 287680 443642 287736
rect 443698 287680 443703 287736
rect 267660 287678 443703 287680
rect 267660 287676 267666 287678
rect 443637 287675 443703 287678
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3233 110666 3299 110669
rect -960 110664 3299 110666
rect -960 110608 3238 110664
rect 3294 110608 3299 110664
rect -960 110606 3299 110608
rect -960 110516 480 110606
rect 3233 110603 3299 110606
rect 579705 99514 579771 99517
rect 583520 99514 584960 99604
rect 579705 99512 584960 99514
rect 579705 99456 579710 99512
rect 579766 99456 584960 99512
rect 579705 99454 584960 99456
rect 579705 99451 579771 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 579981 86186 580047 86189
rect 583520 86186 584960 86276
rect 579981 86184 584960 86186
rect 579981 86128 579986 86184
rect 580042 86128 584960 86184
rect 579981 86126 584960 86128
rect 579981 86123 580047 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 579797 59666 579863 59669
rect 583520 59666 584960 59756
rect 579797 59664 584960 59666
rect 579797 59608 579802 59664
rect 579858 59608 584960 59664
rect 579797 59606 584960 59608
rect 579797 59603 579863 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 580441 19818 580507 19821
rect 583520 19818 584960 19908
rect 580441 19816 584960 19818
rect 580441 19760 580446 19816
rect 580502 19760 584960 19816
rect 580441 19758 584960 19760
rect 580441 19755 580507 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect 583520 6476 584960 6566
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 11145 3498 11211 3501
rect 237373 3498 237439 3501
rect 11145 3496 237439 3498
rect 11145 3440 11150 3496
rect 11206 3440 237378 3496
rect 237434 3440 237439 3496
rect 11145 3438 237439 3440
rect 11145 3435 11211 3438
rect 237373 3435 237439 3438
rect 382549 3498 382615 3501
rect 479333 3498 479399 3501
rect 382549 3496 479399 3498
rect 382549 3440 382554 3496
rect 382610 3440 479338 3496
rect 479394 3440 479399 3496
rect 382549 3438 479399 3440
rect 382549 3435 382615 3438
rect 479333 3435 479399 3438
rect 5257 3362 5323 3365
rect 236269 3362 236335 3365
rect 5257 3360 236335 3362
rect 5257 3304 5262 3360
rect 5318 3304 236274 3360
rect 236330 3304 236335 3360
rect 5257 3302 236335 3304
rect 5257 3299 5323 3302
rect 236269 3299 236335 3302
rect 277117 3362 277183 3365
rect 320265 3362 320331 3365
rect 277117 3360 320331 3362
rect 277117 3304 277122 3360
rect 277178 3304 320270 3360
rect 320326 3304 320331 3360
rect 277117 3302 320331 3304
rect 277117 3299 277183 3302
rect 320265 3299 320331 3302
rect 414381 3362 414447 3365
rect 583385 3362 583451 3365
rect 414381 3360 583451 3362
rect 414381 3304 414386 3360
rect 414442 3304 583390 3360
rect 583446 3304 583451 3360
rect 414381 3302 583451 3304
rect 414381 3299 414447 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 402100 459716 402164 459780
rect 237972 457404 238036 457468
rect 240732 457404 240796 457468
rect 242756 457404 242820 457468
rect 244044 457404 244108 457468
rect 246804 457404 246868 457468
rect 248276 457464 248340 457468
rect 248276 457408 248290 457464
rect 248290 457408 248340 457464
rect 248276 457404 248340 457408
rect 251036 457404 251100 457468
rect 252324 457404 252388 457468
rect 253612 457404 253676 457468
rect 256556 457464 256620 457468
rect 256556 457408 256570 457464
rect 256570 457408 256620 457464
rect 256556 457404 256620 457408
rect 257844 457404 257908 457468
rect 259316 457464 259380 457468
rect 259316 457408 259330 457464
rect 259330 457408 259380 457464
rect 259316 457404 259380 457408
rect 262076 457404 262140 457468
rect 263364 457404 263428 457468
rect 264836 457404 264900 457468
rect 266124 457464 266188 457468
rect 266124 457408 266138 457464
rect 266138 457408 266188 457464
rect 266124 457404 266188 457408
rect 267596 457464 267660 457468
rect 267596 457408 267610 457464
rect 267610 457408 267660 457464
rect 267596 457404 267660 457408
rect 268884 457404 268948 457468
rect 271092 457404 271156 457468
rect 273852 457404 273916 457468
rect 383700 457404 383764 457468
rect 384988 457404 385052 457468
rect 387748 457404 387812 457468
rect 389220 457404 389284 457468
rect 393452 457464 393516 457468
rect 393452 457408 393502 457464
rect 393502 457408 393516 457464
rect 393452 457404 393516 457408
rect 394740 457404 394804 457468
rect 396580 457404 396644 457468
rect 398788 457404 398852 457468
rect 400260 457404 400324 457468
rect 403020 457464 403084 457468
rect 403020 457408 403034 457464
rect 403034 457408 403084 457464
rect 403020 457404 403084 457408
rect 404308 457464 404372 457468
rect 404308 457408 404358 457464
rect 404358 457408 404372 457464
rect 404308 457404 404372 457408
rect 405780 457404 405844 457468
rect 408724 457404 408788 457468
rect 409828 457404 409892 457468
rect 411300 457404 411364 457468
rect 400260 337316 400324 337380
rect 384988 336772 385052 336836
rect 405780 334596 405844 334660
rect 409828 333236 409892 333300
rect 251036 331740 251100 331804
rect 259316 330380 259380 330444
rect 264836 329020 264900 329084
rect 268884 327660 268948 327724
rect 237972 326300 238036 326364
rect 271092 324396 271156 324460
rect 242756 323580 242820 323644
rect 246804 322084 246868 322148
rect 383700 320724 383764 320788
rect 387748 319364 387812 319428
rect 393084 318004 393148 318068
rect 396580 316644 396644 316708
rect 403020 315284 403084 315348
rect 402100 313924 402164 313988
rect 273852 311884 273916 311948
rect 411300 311068 411364 311132
rect 252324 309708 252388 309772
rect 256556 308348 256620 308412
rect 262076 306988 262140 307052
rect 266124 304132 266188 304196
rect 240732 302772 240796 302836
rect 244044 301412 244108 301476
rect 248276 300052 248340 300116
rect 389220 298692 389284 298756
rect 394740 297332 394804 297396
rect 398788 295972 398852 296036
rect 404308 294476 404372 294540
rect 408724 293116 408788 293180
rect 253612 291756 253676 291820
rect 257844 290396 257908 290460
rect 263364 289036 263428 289100
rect 267596 287676 267660 287740
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 237971 457468 238037 457469
rect 237971 457404 237972 457468
rect 238036 457404 238037 457468
rect 237971 457403 238037 457404
rect 240731 457468 240797 457469
rect 240731 457404 240732 457468
rect 240796 457404 240797 457468
rect 240731 457403 240797 457404
rect 242755 457468 242821 457469
rect 242755 457404 242756 457468
rect 242820 457404 242821 457468
rect 242755 457403 242821 457404
rect 244043 457468 244109 457469
rect 244043 457404 244044 457468
rect 244108 457404 244109 457468
rect 244043 457403 244109 457404
rect 246803 457468 246869 457469
rect 246803 457404 246804 457468
rect 246868 457404 246869 457468
rect 246803 457403 246869 457404
rect 248275 457468 248341 457469
rect 248275 457404 248276 457468
rect 248340 457404 248341 457468
rect 248275 457403 248341 457404
rect 251035 457468 251101 457469
rect 251035 457404 251036 457468
rect 251100 457404 251101 457468
rect 251035 457403 251101 457404
rect 252323 457468 252389 457469
rect 252323 457404 252324 457468
rect 252388 457404 252389 457468
rect 252323 457403 252389 457404
rect 253611 457468 253677 457469
rect 253611 457404 253612 457468
rect 253676 457404 253677 457468
rect 253611 457403 253677 457404
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 237974 326365 238034 457403
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 237971 326364 238037 326365
rect 237971 326300 237972 326364
rect 238036 326300 238037 326364
rect 237971 326299 238037 326300
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 240734 302837 240794 457403
rect 242758 323645 242818 457403
rect 242755 323644 242821 323645
rect 242755 323580 242756 323644
rect 242820 323580 242821 323644
rect 242755 323579 242821 323580
rect 240731 302836 240797 302837
rect 240731 302772 240732 302836
rect 240796 302772 240797 302836
rect 240731 302771 240797 302772
rect 244046 301477 244106 457403
rect 246806 322149 246866 457403
rect 246803 322148 246869 322149
rect 246803 322084 246804 322148
rect 246868 322084 246869 322148
rect 246803 322083 246869 322084
rect 244043 301476 244109 301477
rect 244043 301412 244044 301476
rect 244108 301412 244109 301476
rect 244043 301411 244109 301412
rect 248278 300117 248338 457403
rect 251038 331805 251098 457403
rect 251035 331804 251101 331805
rect 251035 331740 251036 331804
rect 251100 331740 251101 331804
rect 251035 331739 251101 331740
rect 252326 309773 252386 457403
rect 252323 309772 252389 309773
rect 252323 309708 252324 309772
rect 252388 309708 252389 309772
rect 252323 309707 252389 309708
rect 248275 300116 248341 300117
rect 248275 300052 248276 300116
rect 248340 300052 248341 300116
rect 248275 300051 248341 300052
rect 253614 291821 253674 457403
rect 253794 435454 254414 470898
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 256555 457468 256621 457469
rect 256555 457404 256556 457468
rect 256620 457404 256621 457468
rect 256555 457403 256621 457404
rect 257843 457468 257909 457469
rect 257843 457404 257844 457468
rect 257908 457404 257909 457468
rect 257843 457403 257909 457404
rect 259315 457468 259381 457469
rect 259315 457404 259316 457468
rect 259380 457404 259381 457468
rect 259315 457403 259381 457404
rect 262075 457468 262141 457469
rect 262075 457404 262076 457468
rect 262140 457404 262141 457468
rect 262075 457403 262141 457404
rect 263363 457468 263429 457469
rect 263363 457404 263364 457468
rect 263428 457404 263429 457468
rect 263363 457403 263429 457404
rect 264835 457468 264901 457469
rect 264835 457404 264836 457468
rect 264900 457404 264901 457468
rect 264835 457403 264901 457404
rect 266123 457468 266189 457469
rect 266123 457404 266124 457468
rect 266188 457404 266189 457468
rect 266123 457403 266189 457404
rect 267595 457468 267661 457469
rect 267595 457404 267596 457468
rect 267660 457404 267661 457468
rect 267595 457403 267661 457404
rect 268883 457468 268949 457469
rect 268883 457404 268884 457468
rect 268948 457404 268949 457468
rect 268883 457403 268949 457404
rect 271091 457468 271157 457469
rect 271091 457404 271092 457468
rect 271156 457404 271157 457468
rect 271091 457403 271157 457404
rect 254568 453454 254888 453486
rect 254568 453218 254610 453454
rect 254846 453218 254888 453454
rect 254568 453134 254888 453218
rect 254568 452898 254610 453134
rect 254846 452898 254888 453134
rect 254568 452866 254888 452898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 254568 417454 254888 417486
rect 254568 417218 254610 417454
rect 254846 417218 254888 417454
rect 254568 417134 254888 417218
rect 254568 416898 254610 417134
rect 254846 416898 254888 417134
rect 254568 416866 254888 416898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253611 291820 253677 291821
rect 253611 291756 253612 291820
rect 253676 291756 253677 291820
rect 253611 291755 253677 291756
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 253794 291454 254414 326898
rect 256558 308413 256618 457403
rect 256555 308412 256621 308413
rect 256555 308348 256556 308412
rect 256620 308348 256621 308412
rect 256555 308347 256621 308348
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 257846 290461 257906 457403
rect 259318 330445 259378 457403
rect 259315 330444 259381 330445
rect 259315 330380 259316 330444
rect 259380 330380 259381 330444
rect 259315 330379 259381 330380
rect 262078 307053 262138 457403
rect 262075 307052 262141 307053
rect 262075 306988 262076 307052
rect 262140 306988 262141 307052
rect 262075 306987 262141 306988
rect 257843 290460 257909 290461
rect 257843 290396 257844 290460
rect 257908 290396 257909 290460
rect 257843 290395 257909 290396
rect 263366 289101 263426 457403
rect 264838 329085 264898 457403
rect 264835 329084 264901 329085
rect 264835 329020 264836 329084
rect 264900 329020 264901 329084
rect 264835 329019 264901 329020
rect 266126 304197 266186 457403
rect 266123 304196 266189 304197
rect 266123 304132 266124 304196
rect 266188 304132 266189 304196
rect 266123 304131 266189 304132
rect 263363 289100 263429 289101
rect 263363 289036 263364 289100
rect 263428 289036 263429 289100
rect 263363 289035 263429 289036
rect 267598 287741 267658 457403
rect 268886 327725 268946 457403
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 268883 327724 268949 327725
rect 268883 327660 268884 327724
rect 268948 327660 268949 327724
rect 268883 327659 268949 327660
rect 271094 324461 271154 457403
rect 271794 453454 272414 488898
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 273851 457468 273917 457469
rect 273851 457404 273852 457468
rect 273916 457404 273917 457468
rect 273851 457403 273917 457404
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271091 324460 271157 324461
rect 271091 324396 271092 324460
rect 271156 324396 271157 324460
rect 271091 324395 271157 324396
rect 271794 309454 272414 344898
rect 273854 311949 273914 457403
rect 285288 453454 285608 453486
rect 285288 453218 285330 453454
rect 285566 453218 285608 453454
rect 285288 453134 285608 453218
rect 285288 452898 285330 453134
rect 285566 452898 285608 453134
rect 285288 452866 285608 452898
rect 289794 435454 290414 470898
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 285288 417454 285608 417486
rect 285288 417218 285330 417454
rect 285566 417218 285608 417454
rect 285288 417134 285608 417218
rect 285288 416898 285330 417134
rect 285566 416898 285608 417134
rect 285288 416866 285608 416898
rect 289794 399454 290414 434898
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 307794 417454 308414 452898
rect 316008 453454 316328 453486
rect 316008 453218 316050 453454
rect 316286 453218 316328 453454
rect 316008 453134 316328 453218
rect 316008 452898 316050 453134
rect 316286 452898 316328 453134
rect 316008 452866 316328 452898
rect 325794 435454 326414 470898
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 285288 381454 285608 381486
rect 285288 381218 285330 381454
rect 285566 381218 285608 381454
rect 285288 381134 285608 381218
rect 285288 380898 285330 381134
rect 285566 380898 285608 381134
rect 285288 380866 285608 380898
rect 289794 363454 290414 398898
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 307794 381454 308414 416898
rect 316008 417454 316328 417486
rect 316008 417218 316050 417454
rect 316286 417218 316328 417454
rect 316008 417134 316328 417218
rect 316008 416898 316050 417134
rect 316286 416898 316328 417134
rect 316008 416866 316328 416898
rect 325794 399454 326414 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 343794 417454 344414 452898
rect 346728 453454 347048 453486
rect 346728 453218 346770 453454
rect 347006 453218 347048 453454
rect 346728 453134 347048 453218
rect 346728 452898 346770 453134
rect 347006 452898 347048 453134
rect 346728 452866 347048 452898
rect 361794 435454 362414 470898
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 377448 453454 377768 453486
rect 377448 453218 377490 453454
rect 377726 453218 377768 453454
rect 377448 453134 377768 453218
rect 377448 452898 377490 453134
rect 377726 452898 377768 453134
rect 377448 452866 377768 452898
rect 379794 453454 380414 488898
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 383699 457468 383765 457469
rect 383699 457404 383700 457468
rect 383764 457404 383765 457468
rect 383699 457403 383765 457404
rect 384987 457468 385053 457469
rect 384987 457404 384988 457468
rect 385052 457404 385053 457468
rect 384987 457403 385053 457404
rect 387747 457468 387813 457469
rect 387747 457404 387748 457468
rect 387812 457404 387813 457468
rect 387747 457403 387813 457404
rect 389219 457468 389285 457469
rect 389219 457404 389220 457468
rect 389284 457404 389285 457468
rect 389219 457403 389285 457404
rect 393451 457468 393517 457469
rect 393451 457404 393452 457468
rect 393516 457404 393517 457468
rect 393451 457403 393517 457404
rect 394739 457468 394805 457469
rect 394739 457404 394740 457468
rect 394804 457404 394805 457468
rect 394739 457403 394805 457404
rect 396579 457468 396645 457469
rect 396579 457404 396580 457468
rect 396644 457404 396645 457468
rect 396579 457403 396645 457404
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 361794 435218 361826 435454
rect 362062 435218 362130 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362130 435134
rect 362382 434898 362414 435134
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 289794 327454 290414 362898
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 273851 311948 273917 311949
rect 273851 311884 273852 311948
rect 273916 311884 273917 311948
rect 273851 311883 273917 311884
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 267595 287740 267661 287741
rect 267595 287676 267596 287740
rect 267660 287676 267661 287740
rect 267595 287675 267661 287676
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 307794 345454 308414 380898
rect 316008 381454 316328 381486
rect 316008 381218 316050 381454
rect 316286 381218 316328 381454
rect 316008 381134 316328 381218
rect 316008 380898 316050 381134
rect 316286 380898 316328 381134
rect 316008 380866 316328 380898
rect 325794 363454 326414 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 343794 381454 344414 416898
rect 346728 417454 347048 417486
rect 346728 417218 346770 417454
rect 347006 417218 347048 417454
rect 346728 417134 347048 417218
rect 346728 416898 346770 417134
rect 347006 416898 347048 417134
rect 346728 416866 347048 416898
rect 361794 399454 362414 434898
rect 377448 417454 377768 417486
rect 377448 417218 377490 417454
rect 377726 417218 377768 417454
rect 377448 417134 377768 417218
rect 377448 416898 377490 417134
rect 377726 416898 377768 417134
rect 377448 416866 377768 416898
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 361794 399218 361826 399454
rect 362062 399218 362130 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362130 399134
rect 362382 398898 362414 399134
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 316008 345454 316328 345486
rect 316008 345218 316050 345454
rect 316286 345218 316328 345454
rect 316008 345134 316328 345218
rect 316008 344898 316050 345134
rect 316286 344898 316328 345134
rect 316008 344866 316328 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 325794 327454 326414 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 343794 345454 344414 380898
rect 346728 381454 347048 381486
rect 346728 381218 346770 381454
rect 347006 381218 347048 381454
rect 346728 381134 347048 381218
rect 346728 380898 346770 381134
rect 347006 380898 347048 381134
rect 346728 380866 347048 380898
rect 361794 363454 362414 398898
rect 377448 381454 377768 381486
rect 377448 381218 377490 381454
rect 377726 381218 377768 381454
rect 377448 381134 377768 381218
rect 377448 380898 377490 381134
rect 377726 380898 377768 381134
rect 377448 380866 377768 380898
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 361794 363218 361826 363454
rect 362062 363218 362130 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362130 363134
rect 362382 362898 362414 363134
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 346728 345454 347048 345486
rect 346728 345218 346770 345454
rect 347006 345218 347048 345454
rect 346728 345134 347048 345218
rect 346728 344898 346770 345134
rect 347006 344898 347048 345134
rect 346728 344866 347048 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 361794 327454 362414 362898
rect 377448 345454 377768 345486
rect 377448 345218 377490 345454
rect 377726 345218 377768 345454
rect 377448 345134 377768 345218
rect 377448 344898 377490 345134
rect 377726 344898 377768 345134
rect 377448 344866 377768 344898
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 379794 309454 380414 344898
rect 383702 320789 383762 457403
rect 384990 336837 385050 457403
rect 384987 336836 385053 336837
rect 384987 336772 384988 336836
rect 385052 336772 385053 336836
rect 384987 336771 385053 336772
rect 383699 320788 383765 320789
rect 383699 320724 383700 320788
rect 383764 320724 383765 320788
rect 383699 320723 383765 320724
rect 387750 319429 387810 457403
rect 387747 319428 387813 319429
rect 387747 319364 387748 319428
rect 387812 319364 387813 319428
rect 387747 319363 387813 319364
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 389222 298757 389282 457403
rect 392808 435454 393128 435486
rect 392808 435218 392850 435454
rect 393086 435218 393128 435454
rect 392808 435134 393128 435218
rect 392808 434898 392850 435134
rect 393086 434898 393128 435134
rect 392808 434866 393128 434898
rect 392808 399454 393128 399486
rect 392808 399218 392850 399454
rect 393086 399218 393128 399454
rect 392808 399134 393128 399218
rect 392808 398898 392850 399134
rect 393086 398898 393128 399134
rect 392808 398866 393128 398898
rect 392808 363454 393128 363486
rect 392808 363218 392850 363454
rect 393086 363218 393128 363454
rect 392808 363134 393128 363218
rect 392808 362898 392850 363134
rect 393086 362898 393128 363134
rect 392808 362866 393128 362898
rect 393454 339690 393514 457403
rect 393086 339630 393514 339690
rect 393086 318069 393146 339630
rect 393083 318068 393149 318069
rect 393083 318004 393084 318068
rect 393148 318004 393149 318068
rect 393083 318003 393149 318004
rect 389219 298756 389285 298757
rect 389219 298692 389220 298756
rect 389284 298692 389285 298756
rect 389219 298691 389285 298692
rect 394742 297397 394802 457403
rect 396582 316709 396642 457403
rect 397794 435454 398414 470898
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 402099 459780 402165 459781
rect 402099 459716 402100 459780
rect 402164 459716 402165 459780
rect 402099 459715 402165 459716
rect 398787 457468 398853 457469
rect 398787 457404 398788 457468
rect 398852 457404 398853 457468
rect 398787 457403 398853 457404
rect 400259 457468 400325 457469
rect 400259 457404 400260 457468
rect 400324 457404 400325 457468
rect 400259 457403 400325 457404
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 398790 331230 398850 457403
rect 400262 337381 400322 457403
rect 400259 337380 400325 337381
rect 400259 337316 400260 337380
rect 400324 337316 400325 337380
rect 400259 337315 400325 337316
rect 398790 331170 399034 331230
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 396579 316708 396645 316709
rect 396579 316644 396580 316708
rect 396644 316644 396645 316708
rect 396579 316643 396645 316644
rect 394739 297396 394805 297397
rect 394739 297332 394740 297396
rect 394804 297332 394805 297396
rect 394739 297331 394805 297332
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 397794 291454 398414 326898
rect 398974 321570 399034 331170
rect 398790 321510 399034 321570
rect 398790 296037 398850 321510
rect 402102 313989 402162 459715
rect 403019 457468 403085 457469
rect 403019 457404 403020 457468
rect 403084 457404 403085 457468
rect 403019 457403 403085 457404
rect 404307 457468 404373 457469
rect 404307 457404 404308 457468
rect 404372 457404 404373 457468
rect 404307 457403 404373 457404
rect 405779 457468 405845 457469
rect 405779 457404 405780 457468
rect 405844 457404 405845 457468
rect 405779 457403 405845 457404
rect 408723 457468 408789 457469
rect 408723 457404 408724 457468
rect 408788 457404 408789 457468
rect 408723 457403 408789 457404
rect 409827 457468 409893 457469
rect 409827 457404 409828 457468
rect 409892 457404 409893 457468
rect 409827 457403 409893 457404
rect 411299 457468 411365 457469
rect 411299 457404 411300 457468
rect 411364 457404 411365 457468
rect 411299 457403 411365 457404
rect 403022 315349 403082 457403
rect 403019 315348 403085 315349
rect 403019 315284 403020 315348
rect 403084 315284 403085 315348
rect 403019 315283 403085 315284
rect 402099 313988 402165 313989
rect 402099 313924 402100 313988
rect 402164 313924 402165 313988
rect 402099 313923 402165 313924
rect 398787 296036 398853 296037
rect 398787 295972 398788 296036
rect 398852 295972 398853 296036
rect 398787 295971 398853 295972
rect 404310 294541 404370 457403
rect 405782 334661 405842 457403
rect 408168 453454 408488 453486
rect 408168 453218 408210 453454
rect 408446 453218 408488 453454
rect 408168 453134 408488 453218
rect 408168 452898 408210 453134
rect 408446 452898 408488 453134
rect 408168 452866 408488 452898
rect 408168 417454 408488 417486
rect 408168 417218 408210 417454
rect 408446 417218 408488 417454
rect 408168 417134 408488 417218
rect 408168 416898 408210 417134
rect 408446 416898 408488 417134
rect 408168 416866 408488 416898
rect 408168 381454 408488 381486
rect 408168 381218 408210 381454
rect 408446 381218 408488 381454
rect 408168 381134 408488 381218
rect 408168 380898 408210 381134
rect 408446 380898 408488 381134
rect 408168 380866 408488 380898
rect 408168 345454 408488 345486
rect 408168 345218 408210 345454
rect 408446 345218 408488 345454
rect 408168 345134 408488 345218
rect 408168 344898 408210 345134
rect 408446 344898 408488 345134
rect 408168 344866 408488 344898
rect 405779 334660 405845 334661
rect 405779 334596 405780 334660
rect 405844 334596 405845 334660
rect 405779 334595 405845 334596
rect 404307 294540 404373 294541
rect 404307 294476 404308 294540
rect 404372 294476 404373 294540
rect 404307 294475 404373 294476
rect 408726 293181 408786 457403
rect 409830 333301 409890 457403
rect 409827 333300 409893 333301
rect 409827 333236 409828 333300
rect 409892 333236 409893 333300
rect 409827 333235 409893 333236
rect 411302 311133 411362 457403
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 411299 311132 411365 311133
rect 411299 311068 411300 311132
rect 411364 311068 411365 311132
rect 411299 311067 411365 311068
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 408723 293180 408789 293181
rect 408723 293116 408724 293180
rect 408788 293116 408789 293180
rect 408723 293115 408789 293116
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 577794 704838 578414 705830
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 254610 453218 254846 453454
rect 254610 452898 254846 453134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 254610 417218 254846 417454
rect 254610 416898 254846 417134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 285330 453218 285566 453454
rect 285330 452898 285566 453134
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 285330 417218 285566 417454
rect 285330 416898 285566 417134
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 316050 453218 316286 453454
rect 316050 452898 316286 453134
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 285330 381218 285566 381454
rect 285330 380898 285566 381134
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 316050 417218 316286 417454
rect 316050 416898 316286 417134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 346770 453218 347006 453454
rect 346770 452898 347006 453134
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 377490 453218 377726 453454
rect 377490 452898 377726 453134
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 361826 435218 362062 435454
rect 362130 435218 362382 435454
rect 361826 434898 362062 435134
rect 362130 434898 362382 435134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 316050 381218 316286 381454
rect 316050 380898 316286 381134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 346770 417218 347006 417454
rect 346770 416898 347006 417134
rect 377490 417218 377726 417454
rect 377490 416898 377726 417134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 361826 399218 362062 399454
rect 362130 399218 362382 399454
rect 361826 398898 362062 399134
rect 362130 398898 362382 399134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 316050 345218 316286 345454
rect 316050 344898 316286 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 346770 381218 347006 381454
rect 346770 380898 347006 381134
rect 377490 381218 377726 381454
rect 377490 380898 377726 381134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 361826 363218 362062 363454
rect 362130 363218 362382 363454
rect 361826 362898 362062 363134
rect 362130 362898 362382 363134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 346770 345218 347006 345454
rect 346770 344898 347006 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 377490 345218 377726 345454
rect 377490 344898 377726 345134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 392850 435218 393086 435454
rect 392850 434898 393086 435134
rect 392850 399218 393086 399454
rect 392850 398898 393086 399134
rect 392850 363218 393086 363454
rect 392850 362898 393086 363134
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 408210 453218 408446 453454
rect 408210 452898 408446 453134
rect 408210 417218 408446 417454
rect 408210 416898 408446 417134
rect 408210 381218 408446 381454
rect 408210 380898 408446 381134
rect 408210 345218 408446 345454
rect 408210 344898 408446 345134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 254610 453454
rect 254846 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 285330 453454
rect 285566 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 316050 453454
rect 316286 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 346770 453454
rect 347006 453218 377490 453454
rect 377726 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 408210 453454
rect 408446 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 254610 453134
rect 254846 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 285330 453134
rect 285566 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 316050 453134
rect 316286 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 346770 453134
rect 347006 452898 377490 453134
rect 377726 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 408210 453134
rect 408446 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 239250 435454
rect 239486 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 269970 435454
rect 270206 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 300690 435454
rect 300926 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 331410 435454
rect 331646 435218 361826 435454
rect 362062 435218 362130 435454
rect 362382 435218 392850 435454
rect 393086 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 239250 435134
rect 239486 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 269970 435134
rect 270206 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 300690 435134
rect 300926 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 331410 435134
rect 331646 434898 361826 435134
rect 362062 434898 362130 435134
rect 362382 434898 392850 435134
rect 393086 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 254610 417454
rect 254846 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 285330 417454
rect 285566 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 316050 417454
rect 316286 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 346770 417454
rect 347006 417218 377490 417454
rect 377726 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 408210 417454
rect 408446 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 254610 417134
rect 254846 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 285330 417134
rect 285566 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 316050 417134
rect 316286 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 346770 417134
rect 347006 416898 377490 417134
rect 377726 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 408210 417134
rect 408446 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 239250 399454
rect 239486 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 269970 399454
rect 270206 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 300690 399454
rect 300926 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 331410 399454
rect 331646 399218 361826 399454
rect 362062 399218 362130 399454
rect 362382 399218 392850 399454
rect 393086 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 239250 399134
rect 239486 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 269970 399134
rect 270206 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 300690 399134
rect 300926 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 331410 399134
rect 331646 398898 361826 399134
rect 362062 398898 362130 399134
rect 362382 398898 392850 399134
rect 393086 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 254610 381454
rect 254846 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 285330 381454
rect 285566 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 316050 381454
rect 316286 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 346770 381454
rect 347006 381218 377490 381454
rect 377726 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 408210 381454
rect 408446 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 254610 381134
rect 254846 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 285330 381134
rect 285566 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 316050 381134
rect 316286 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 346770 381134
rect 347006 380898 377490 381134
rect 377726 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 408210 381134
rect 408446 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 239250 363454
rect 239486 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 269970 363454
rect 270206 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 300690 363454
rect 300926 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 331410 363454
rect 331646 363218 361826 363454
rect 362062 363218 362130 363454
rect 362382 363218 392850 363454
rect 393086 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 239250 363134
rect 239486 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 269970 363134
rect 270206 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 300690 363134
rect 300926 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 331410 363134
rect 331646 362898 361826 363134
rect 362062 362898 362130 363134
rect 362382 362898 392850 363134
rect 393086 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 254610 345454
rect 254846 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 285330 345454
rect 285566 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 316050 345454
rect 316286 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 346770 345454
rect 347006 345218 377490 345454
rect 377726 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 408210 345454
rect 408446 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 254610 345134
rect 254846 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 285330 345134
rect 285566 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 316050 345134
rect 316286 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 346770 345134
rect 347006 344898 377490 345134
rect 377726 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 408210 345134
rect 408446 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use user_proj_example  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box 105 0 179846 120000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 532 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 532 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 532 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 532 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 533 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 535 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 536 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 537 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 538 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 539 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 540 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 541 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 542 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 543 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 544 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 545 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 546 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 547 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 548 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 549 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 550 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 551 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 552 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 553 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 554 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 555 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 556 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 557 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 558 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 559 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 560 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 561 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 562 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 563 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 564 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 565 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 566 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 567 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 568 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 569 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 570 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 571 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 572 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 573 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 574 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 575 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 576 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 577 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 578 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 579 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 580 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 581 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 582 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 583 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 584 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 585 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 586 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 587 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 588 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 589 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 590 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 591 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 592 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 593 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 594 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 595 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 596 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 597 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 598 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 599 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 600 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 601 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 602 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 603 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 604 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 605 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 606 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 607 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 608 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 609 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 610 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 611 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 612 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 613 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 614 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 615 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 616 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 617 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 618 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 619 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 620 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 621 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 622 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 623 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 624 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 625 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 626 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 627 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 628 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 629 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 630 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 631 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 632 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 633 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 634 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 635 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 636 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 637 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
